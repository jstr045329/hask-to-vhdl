library IEEE;
use IEEE.std_logic_1164.ALL;
use IEEE.numeric_std.ALL;


entity ArbSetLowLayerNode is
    port (
        clk : in std_logic;
        rst : in std_logic
    );
end ArbSetLowLayerNode;


architecture behavioral_ArbSetLowLayerNode of ArbSetLowLayerNode is
begin


end behavioral_ArbSetLowLayerNode;

