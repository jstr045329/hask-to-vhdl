library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.PrefixFunctions.all;


package SingleCyclePipelinedFunctions is


function large_and (
    x_000000_000000 : std_logic;
    x_000001_000000 : std_logic := '0';
    x_000002_000000 : std_logic := '0';
    x_000003_000000 : std_logic := '0';
    x_000004_000000 : std_logic := '0';
    x_000005_000000 : std_logic := '0';
    x_000006_000000 : std_logic := '0';
    x_000007_000000 : std_logic := '0';
    x_000008_000000 : std_logic := '0';
    x_000009_000000 : std_logic := '0';
    x_000010_000000 : std_logic := '0';
    x_000011_000000 : std_logic := '0';
    x_000012_000000 : std_logic := '0';
    x_000013_000000 : std_logic := '0';
    x_000014_000000 : std_logic := '0';
    x_000015_000000 : std_logic := '0';
    x_000016_000000 : std_logic := '0';
    x_000017_000000 : std_logic := '0';
    x_000018_000000 : std_logic := '0';
    x_000019_000000 : std_logic := '0';
    x_000020_000000 : std_logic := '0';
    x_000021_000000 : std_logic := '0';
    x_000022_000000 : std_logic := '0';
    x_000023_000000 : std_logic := '0';
    x_000024_000000 : std_logic := '0';
    x_000025_000000 : std_logic := '0';
    x_000026_000000 : std_logic := '0';
    x_000027_000000 : std_logic := '0';
    x_000028_000000 : std_logic := '0';
    x_000029_000000 : std_logic := '0';
    x_000030_000000 : std_logic := '0';
    x_000031_000000 : std_logic := '0';
    x_000032_000000 : std_logic := '0';
    x_000033_000000 : std_logic := '0';
    x_000034_000000 : std_logic := '0';
    x_000035_000000 : std_logic := '0';
    x_000036_000000 : std_logic := '0';
    x_000037_000000 : std_logic := '0';
    x_000038_000000 : std_logic := '0';
    x_000039_000000 : std_logic := '0';
    x_000040_000000 : std_logic := '0';
    x_000041_000000 : std_logic := '0';
    x_000042_000000 : std_logic := '0';
    x_000043_000000 : std_logic := '0';
    x_000044_000000 : std_logic := '0';
    x_000045_000000 : std_logic := '0';
    x_000046_000000 : std_logic := '0';
    x_000047_000000 : std_logic := '0';
    x_000048_000000 : std_logic := '0';
    x_000049_000000 : std_logic := '0';
    x_000050_000000 : std_logic := '0';
    x_000051_000000 : std_logic := '0';
    x_000052_000000 : std_logic := '0';
    x_000053_000000 : std_logic := '0';
    x_000054_000000 : std_logic := '0';
    x_000055_000000 : std_logic := '0';
    x_000056_000000 : std_logic := '0';
    x_000057_000000 : std_logic := '0';
    x_000058_000000 : std_logic := '0';
    x_000059_000000 : std_logic := '0';
    x_000060_000000 : std_logic := '0';
    x_000061_000000 : std_logic := '0';
    x_000062_000000 : std_logic := '0';
    x_000063_000000 : std_logic := '0';
    x_000064_000000 : std_logic := '0';
    x_000065_000000 : std_logic := '0';
    x_000066_000000 : std_logic := '0';
    x_000067_000000 : std_logic := '0';
    x_000068_000000 : std_logic := '0';
    x_000069_000000 : std_logic := '0';
    x_000070_000000 : std_logic := '0';
    x_000071_000000 : std_logic := '0';
    x_000072_000000 : std_logic := '0';
    x_000073_000000 : std_logic := '0';
    x_000074_000000 : std_logic := '0';
    x_000075_000000 : std_logic := '0';
    x_000076_000000 : std_logic := '0';
    x_000077_000000 : std_logic := '0';
    x_000078_000000 : std_logic := '0';
    x_000079_000000 : std_logic := '0';
    x_000080_000000 : std_logic := '0';
    x_000081_000000 : std_logic := '0';
    x_000082_000000 : std_logic := '0';
    x_000083_000000 : std_logic := '0';
    x_000084_000000 : std_logic := '0';
    x_000085_000000 : std_logic := '0';
    x_000086_000000 : std_logic := '0';
    x_000087_000000 : std_logic := '0';
    x_000088_000000 : std_logic := '0';
    x_000089_000000 : std_logic := '0';
    x_000090_000000 : std_logic := '0';
    x_000091_000000 : std_logic := '0';
    x_000092_000000 : std_logic := '0';
    x_000093_000000 : std_logic := '0';
    x_000094_000000 : std_logic := '0';
    x_000095_000000 : std_logic := '0';
    x_000096_000000 : std_logic := '0';
    x_000097_000000 : std_logic := '0';
    x_000098_000000 : std_logic := '0';
    x_000099_000000 : std_logic := '0';
    x_000100_000000 : std_logic := '0';
    x_000101_000000 : std_logic := '0';
    x_000102_000000 : std_logic := '0';
    x_000103_000000 : std_logic := '0';
    x_000104_000000 : std_logic := '0';
    x_000105_000000 : std_logic := '0';
    x_000106_000000 : std_logic := '0';
    x_000107_000000 : std_logic := '0';
    x_000108_000000 : std_logic := '0';
    x_000109_000000 : std_logic := '0';
    x_000110_000000 : std_logic := '0';
    x_000111_000000 : std_logic := '0';
    x_000112_000000 : std_logic := '0';
    x_000113_000000 : std_logic := '0';
    x_000114_000000 : std_logic := '0';
    x_000115_000000 : std_logic := '0';
    x_000116_000000 : std_logic := '0';
    x_000117_000000 : std_logic := '0';
    x_000118_000000 : std_logic := '0';
    x_000119_000000 : std_logic := '0';
    x_000120_000000 : std_logic := '0';
    x_000121_000000 : std_logic := '0';
    x_000122_000000 : std_logic := '0';
    x_000123_000000 : std_logic := '0';
    x_000124_000000 : std_logic := '0';
    x_000125_000000 : std_logic := '0';
    x_000126_000000 : std_logic := '0';
    x_000127_000000 : std_logic := '0') return std_logic;
    

function large_or (
    x_000000_000000 : std_logic;
    x_000001_000000 : std_logic := '0';
    x_000002_000000 : std_logic := '0';
    x_000003_000000 : std_logic := '0';
    x_000004_000000 : std_logic := '0';
    x_000005_000000 : std_logic := '0';
    x_000006_000000 : std_logic := '0';
    x_000007_000000 : std_logic := '0';
    x_000008_000000 : std_logic := '0';
    x_000009_000000 : std_logic := '0';
    x_000010_000000 : std_logic := '0';
    x_000011_000000 : std_logic := '0';
    x_000012_000000 : std_logic := '0';
    x_000013_000000 : std_logic := '0';
    x_000014_000000 : std_logic := '0';
    x_000015_000000 : std_logic := '0';
    x_000016_000000 : std_logic := '0';
    x_000017_000000 : std_logic := '0';
    x_000018_000000 : std_logic := '0';
    x_000019_000000 : std_logic := '0';
    x_000020_000000 : std_logic := '0';
    x_000021_000000 : std_logic := '0';
    x_000022_000000 : std_logic := '0';
    x_000023_000000 : std_logic := '0';
    x_000024_000000 : std_logic := '0';
    x_000025_000000 : std_logic := '0';
    x_000026_000000 : std_logic := '0';
    x_000027_000000 : std_logic := '0';
    x_000028_000000 : std_logic := '0';
    x_000029_000000 : std_logic := '0';
    x_000030_000000 : std_logic := '0';
    x_000031_000000 : std_logic := '0';
    x_000032_000000 : std_logic := '0';
    x_000033_000000 : std_logic := '0';
    x_000034_000000 : std_logic := '0';
    x_000035_000000 : std_logic := '0';
    x_000036_000000 : std_logic := '0';
    x_000037_000000 : std_logic := '0';
    x_000038_000000 : std_logic := '0';
    x_000039_000000 : std_logic := '0';
    x_000040_000000 : std_logic := '0';
    x_000041_000000 : std_logic := '0';
    x_000042_000000 : std_logic := '0';
    x_000043_000000 : std_logic := '0';
    x_000044_000000 : std_logic := '0';
    x_000045_000000 : std_logic := '0';
    x_000046_000000 : std_logic := '0';
    x_000047_000000 : std_logic := '0';
    x_000048_000000 : std_logic := '0';
    x_000049_000000 : std_logic := '0';
    x_000050_000000 : std_logic := '0';
    x_000051_000000 : std_logic := '0';
    x_000052_000000 : std_logic := '0';
    x_000053_000000 : std_logic := '0';
    x_000054_000000 : std_logic := '0';
    x_000055_000000 : std_logic := '0';
    x_000056_000000 : std_logic := '0';
    x_000057_000000 : std_logic := '0';
    x_000058_000000 : std_logic := '0';
    x_000059_000000 : std_logic := '0';
    x_000060_000000 : std_logic := '0';
    x_000061_000000 : std_logic := '0';
    x_000062_000000 : std_logic := '0';
    x_000063_000000 : std_logic := '0';
    x_000064_000000 : std_logic := '0';
    x_000065_000000 : std_logic := '0';
    x_000066_000000 : std_logic := '0';
    x_000067_000000 : std_logic := '0';
    x_000068_000000 : std_logic := '0';
    x_000069_000000 : std_logic := '0';
    x_000070_000000 : std_logic := '0';
    x_000071_000000 : std_logic := '0';
    x_000072_000000 : std_logic := '0';
    x_000073_000000 : std_logic := '0';
    x_000074_000000 : std_logic := '0';
    x_000075_000000 : std_logic := '0';
    x_000076_000000 : std_logic := '0';
    x_000077_000000 : std_logic := '0';
    x_000078_000000 : std_logic := '0';
    x_000079_000000 : std_logic := '0';
    x_000080_000000 : std_logic := '0';
    x_000081_000000 : std_logic := '0';
    x_000082_000000 : std_logic := '0';
    x_000083_000000 : std_logic := '0';
    x_000084_000000 : std_logic := '0';
    x_000085_000000 : std_logic := '0';
    x_000086_000000 : std_logic := '0';
    x_000087_000000 : std_logic := '0';
    x_000088_000000 : std_logic := '0';
    x_000089_000000 : std_logic := '0';
    x_000090_000000 : std_logic := '0';
    x_000091_000000 : std_logic := '0';
    x_000092_000000 : std_logic := '0';
    x_000093_000000 : std_logic := '0';
    x_000094_000000 : std_logic := '0';
    x_000095_000000 : std_logic := '0';
    x_000096_000000 : std_logic := '0';
    x_000097_000000 : std_logic := '0';
    x_000098_000000 : std_logic := '0';
    x_000099_000000 : std_logic := '0';
    x_000100_000000 : std_logic := '0';
    x_000101_000000 : std_logic := '0';
    x_000102_000000 : std_logic := '0';
    x_000103_000000 : std_logic := '0';
    x_000104_000000 : std_logic := '0';
    x_000105_000000 : std_logic := '0';
    x_000106_000000 : std_logic := '0';
    x_000107_000000 : std_logic := '0';
    x_000108_000000 : std_logic := '0';
    x_000109_000000 : std_logic := '0';
    x_000110_000000 : std_logic := '0';
    x_000111_000000 : std_logic := '0';
    x_000112_000000 : std_logic := '0';
    x_000113_000000 : std_logic := '0';
    x_000114_000000 : std_logic := '0';
    x_000115_000000 : std_logic := '0';
    x_000116_000000 : std_logic := '0';
    x_000117_000000 : std_logic := '0';
    x_000118_000000 : std_logic := '0';
    x_000119_000000 : std_logic := '0';
    x_000120_000000 : std_logic := '0';
    x_000121_000000 : std_logic := '0';
    x_000122_000000 : std_logic := '0';
    x_000123_000000 : std_logic := '0';
    x_000124_000000 : std_logic := '0';
    x_000125_000000 : std_logic := '0';
    x_000126_000000 : std_logic := '0';
    x_000127_000000 : std_logic := '0') return std_logic;


function large_nand (
    x_000000_000000 : std_logic;
    x_000001_000000 : std_logic := '0';
    x_000002_000000 : std_logic := '0';
    x_000003_000000 : std_logic := '0';
    x_000004_000000 : std_logic := '0';
    x_000005_000000 : std_logic := '0';
    x_000006_000000 : std_logic := '0';
    x_000007_000000 : std_logic := '0';
    x_000008_000000 : std_logic := '0';
    x_000009_000000 : std_logic := '0';
    x_000010_000000 : std_logic := '0';
    x_000011_000000 : std_logic := '0';
    x_000012_000000 : std_logic := '0';
    x_000013_000000 : std_logic := '0';
    x_000014_000000 : std_logic := '0';
    x_000015_000000 : std_logic := '0';
    x_000016_000000 : std_logic := '0';
    x_000017_000000 : std_logic := '0';
    x_000018_000000 : std_logic := '0';
    x_000019_000000 : std_logic := '0';
    x_000020_000000 : std_logic := '0';
    x_000021_000000 : std_logic := '0';
    x_000022_000000 : std_logic := '0';
    x_000023_000000 : std_logic := '0';
    x_000024_000000 : std_logic := '0';
    x_000025_000000 : std_logic := '0';
    x_000026_000000 : std_logic := '0';
    x_000027_000000 : std_logic := '0';
    x_000028_000000 : std_logic := '0';
    x_000029_000000 : std_logic := '0';
    x_000030_000000 : std_logic := '0';
    x_000031_000000 : std_logic := '0';
    x_000032_000000 : std_logic := '0';
    x_000033_000000 : std_logic := '0';
    x_000034_000000 : std_logic := '0';
    x_000035_000000 : std_logic := '0';
    x_000036_000000 : std_logic := '0';
    x_000037_000000 : std_logic := '0';
    x_000038_000000 : std_logic := '0';
    x_000039_000000 : std_logic := '0';
    x_000040_000000 : std_logic := '0';
    x_000041_000000 : std_logic := '0';
    x_000042_000000 : std_logic := '0';
    x_000043_000000 : std_logic := '0';
    x_000044_000000 : std_logic := '0';
    x_000045_000000 : std_logic := '0';
    x_000046_000000 : std_logic := '0';
    x_000047_000000 : std_logic := '0';
    x_000048_000000 : std_logic := '0';
    x_000049_000000 : std_logic := '0';
    x_000050_000000 : std_logic := '0';
    x_000051_000000 : std_logic := '0';
    x_000052_000000 : std_logic := '0';
    x_000053_000000 : std_logic := '0';
    x_000054_000000 : std_logic := '0';
    x_000055_000000 : std_logic := '0';
    x_000056_000000 : std_logic := '0';
    x_000057_000000 : std_logic := '0';
    x_000058_000000 : std_logic := '0';
    x_000059_000000 : std_logic := '0';
    x_000060_000000 : std_logic := '0';
    x_000061_000000 : std_logic := '0';
    x_000062_000000 : std_logic := '0';
    x_000063_000000 : std_logic := '0';
    x_000064_000000 : std_logic := '0';
    x_000065_000000 : std_logic := '0';
    x_000066_000000 : std_logic := '0';
    x_000067_000000 : std_logic := '0';
    x_000068_000000 : std_logic := '0';
    x_000069_000000 : std_logic := '0';
    x_000070_000000 : std_logic := '0';
    x_000071_000000 : std_logic := '0';
    x_000072_000000 : std_logic := '0';
    x_000073_000000 : std_logic := '0';
    x_000074_000000 : std_logic := '0';
    x_000075_000000 : std_logic := '0';
    x_000076_000000 : std_logic := '0';
    x_000077_000000 : std_logic := '0';
    x_000078_000000 : std_logic := '0';
    x_000079_000000 : std_logic := '0';
    x_000080_000000 : std_logic := '0';
    x_000081_000000 : std_logic := '0';
    x_000082_000000 : std_logic := '0';
    x_000083_000000 : std_logic := '0';
    x_000084_000000 : std_logic := '0';
    x_000085_000000 : std_logic := '0';
    x_000086_000000 : std_logic := '0';
    x_000087_000000 : std_logic := '0';
    x_000088_000000 : std_logic := '0';
    x_000089_000000 : std_logic := '0';
    x_000090_000000 : std_logic := '0';
    x_000091_000000 : std_logic := '0';
    x_000092_000000 : std_logic := '0';
    x_000093_000000 : std_logic := '0';
    x_000094_000000 : std_logic := '0';
    x_000095_000000 : std_logic := '0';
    x_000096_000000 : std_logic := '0';
    x_000097_000000 : std_logic := '0';
    x_000098_000000 : std_logic := '0';
    x_000099_000000 : std_logic := '0';
    x_000100_000000 : std_logic := '0';
    x_000101_000000 : std_logic := '0';
    x_000102_000000 : std_logic := '0';
    x_000103_000000 : std_logic := '0';
    x_000104_000000 : std_logic := '0';
    x_000105_000000 : std_logic := '0';
    x_000106_000000 : std_logic := '0';
    x_000107_000000 : std_logic := '0';
    x_000108_000000 : std_logic := '0';
    x_000109_000000 : std_logic := '0';
    x_000110_000000 : std_logic := '0';
    x_000111_000000 : std_logic := '0';
    x_000112_000000 : std_logic := '0';
    x_000113_000000 : std_logic := '0';
    x_000114_000000 : std_logic := '0';
    x_000115_000000 : std_logic := '0';
    x_000116_000000 : std_logic := '0';
    x_000117_000000 : std_logic := '0';
    x_000118_000000 : std_logic := '0';
    x_000119_000000 : std_logic := '0';
    x_000120_000000 : std_logic := '0';
    x_000121_000000 : std_logic := '0';
    x_000122_000000 : std_logic := '0';
    x_000123_000000 : std_logic := '0';
    x_000124_000000 : std_logic := '0';
    x_000125_000000 : std_logic := '0';
    x_000126_000000 : std_logic := '0';
    x_000127_000000 : std_logic := '0') return std_logic;


function large_nor (
    x_000000_000000 : std_logic;
    x_000001_000000 : std_logic := '0';
    x_000002_000000 : std_logic := '0';
    x_000003_000000 : std_logic := '0';
    x_000004_000000 : std_logic := '0';
    x_000005_000000 : std_logic := '0';
    x_000006_000000 : std_logic := '0';
    x_000007_000000 : std_logic := '0';
    x_000008_000000 : std_logic := '0';
    x_000009_000000 : std_logic := '0';
    x_000010_000000 : std_logic := '0';
    x_000011_000000 : std_logic := '0';
    x_000012_000000 : std_logic := '0';
    x_000013_000000 : std_logic := '0';
    x_000014_000000 : std_logic := '0';
    x_000015_000000 : std_logic := '0';
    x_000016_000000 : std_logic := '0';
    x_000017_000000 : std_logic := '0';
    x_000018_000000 : std_logic := '0';
    x_000019_000000 : std_logic := '0';
    x_000020_000000 : std_logic := '0';
    x_000021_000000 : std_logic := '0';
    x_000022_000000 : std_logic := '0';
    x_000023_000000 : std_logic := '0';
    x_000024_000000 : std_logic := '0';
    x_000025_000000 : std_logic := '0';
    x_000026_000000 : std_logic := '0';
    x_000027_000000 : std_logic := '0';
    x_000028_000000 : std_logic := '0';
    x_000029_000000 : std_logic := '0';
    x_000030_000000 : std_logic := '0';
    x_000031_000000 : std_logic := '0';
    x_000032_000000 : std_logic := '0';
    x_000033_000000 : std_logic := '0';
    x_000034_000000 : std_logic := '0';
    x_000035_000000 : std_logic := '0';
    x_000036_000000 : std_logic := '0';
    x_000037_000000 : std_logic := '0';
    x_000038_000000 : std_logic := '0';
    x_000039_000000 : std_logic := '0';
    x_000040_000000 : std_logic := '0';
    x_000041_000000 : std_logic := '0';
    x_000042_000000 : std_logic := '0';
    x_000043_000000 : std_logic := '0';
    x_000044_000000 : std_logic := '0';
    x_000045_000000 : std_logic := '0';
    x_000046_000000 : std_logic := '0';
    x_000047_000000 : std_logic := '0';
    x_000048_000000 : std_logic := '0';
    x_000049_000000 : std_logic := '0';
    x_000050_000000 : std_logic := '0';
    x_000051_000000 : std_logic := '0';
    x_000052_000000 : std_logic := '0';
    x_000053_000000 : std_logic := '0';
    x_000054_000000 : std_logic := '0';
    x_000055_000000 : std_logic := '0';
    x_000056_000000 : std_logic := '0';
    x_000057_000000 : std_logic := '0';
    x_000058_000000 : std_logic := '0';
    x_000059_000000 : std_logic := '0';
    x_000060_000000 : std_logic := '0';
    x_000061_000000 : std_logic := '0';
    x_000062_000000 : std_logic := '0';
    x_000063_000000 : std_logic := '0';
    x_000064_000000 : std_logic := '0';
    x_000065_000000 : std_logic := '0';
    x_000066_000000 : std_logic := '0';
    x_000067_000000 : std_logic := '0';
    x_000068_000000 : std_logic := '0';
    x_000069_000000 : std_logic := '0';
    x_000070_000000 : std_logic := '0';
    x_000071_000000 : std_logic := '0';
    x_000072_000000 : std_logic := '0';
    x_000073_000000 : std_logic := '0';
    x_000074_000000 : std_logic := '0';
    x_000075_000000 : std_logic := '0';
    x_000076_000000 : std_logic := '0';
    x_000077_000000 : std_logic := '0';
    x_000078_000000 : std_logic := '0';
    x_000079_000000 : std_logic := '0';
    x_000080_000000 : std_logic := '0';
    x_000081_000000 : std_logic := '0';
    x_000082_000000 : std_logic := '0';
    x_000083_000000 : std_logic := '0';
    x_000084_000000 : std_logic := '0';
    x_000085_000000 : std_logic := '0';
    x_000086_000000 : std_logic := '0';
    x_000087_000000 : std_logic := '0';
    x_000088_000000 : std_logic := '0';
    x_000089_000000 : std_logic := '0';
    x_000090_000000 : std_logic := '0';
    x_000091_000000 : std_logic := '0';
    x_000092_000000 : std_logic := '0';
    x_000093_000000 : std_logic := '0';
    x_000094_000000 : std_logic := '0';
    x_000095_000000 : std_logic := '0';
    x_000096_000000 : std_logic := '0';
    x_000097_000000 : std_logic := '0';
    x_000098_000000 : std_logic := '0';
    x_000099_000000 : std_logic := '0';
    x_000100_000000 : std_logic := '0';
    x_000101_000000 : std_logic := '0';
    x_000102_000000 : std_logic := '0';
    x_000103_000000 : std_logic := '0';
    x_000104_000000 : std_logic := '0';
    x_000105_000000 : std_logic := '0';
    x_000106_000000 : std_logic := '0';
    x_000107_000000 : std_logic := '0';
    x_000108_000000 : std_logic := '0';
    x_000109_000000 : std_logic := '0';
    x_000110_000000 : std_logic := '0';
    x_000111_000000 : std_logic := '0';
    x_000112_000000 : std_logic := '0';
    x_000113_000000 : std_logic := '0';
    x_000114_000000 : std_logic := '0';
    x_000115_000000 : std_logic := '0';
    x_000116_000000 : std_logic := '0';
    x_000117_000000 : std_logic := '0';
    x_000118_000000 : std_logic := '0';
    x_000119_000000 : std_logic := '0';
    x_000120_000000 : std_logic := '0';
    x_000121_000000 : std_logic := '0';
    x_000122_000000 : std_logic := '0';
    x_000123_000000 : std_logic := '0';
    x_000124_000000 : std_logic := '0';
    x_000125_000000 : std_logic := '0';
    x_000126_000000 : std_logic := '0';
    x_000127_000000 : std_logic := '0') return std_logic;


function large_xor (
    x_000000_000000 : std_logic;
    x_000001_000000 : std_logic := '0';
    x_000002_000000 : std_logic := '0';
    x_000003_000000 : std_logic := '0';
    x_000004_000000 : std_logic := '0';
    x_000005_000000 : std_logic := '0';
    x_000006_000000 : std_logic := '0';
    x_000007_000000 : std_logic := '0';
    x_000008_000000 : std_logic := '0';
    x_000009_000000 : std_logic := '0';
    x_000010_000000 : std_logic := '0';
    x_000011_000000 : std_logic := '0';
    x_000012_000000 : std_logic := '0';
    x_000013_000000 : std_logic := '0';
    x_000014_000000 : std_logic := '0';
    x_000015_000000 : std_logic := '0';
    x_000016_000000 : std_logic := '0';
    x_000017_000000 : std_logic := '0';
    x_000018_000000 : std_logic := '0';
    x_000019_000000 : std_logic := '0';
    x_000020_000000 : std_logic := '0';
    x_000021_000000 : std_logic := '0';
    x_000022_000000 : std_logic := '0';
    x_000023_000000 : std_logic := '0';
    x_000024_000000 : std_logic := '0';
    x_000025_000000 : std_logic := '0';
    x_000026_000000 : std_logic := '0';
    x_000027_000000 : std_logic := '0';
    x_000028_000000 : std_logic := '0';
    x_000029_000000 : std_logic := '0';
    x_000030_000000 : std_logic := '0';
    x_000031_000000 : std_logic := '0';
    x_000032_000000 : std_logic := '0';
    x_000033_000000 : std_logic := '0';
    x_000034_000000 : std_logic := '0';
    x_000035_000000 : std_logic := '0';
    x_000036_000000 : std_logic := '0';
    x_000037_000000 : std_logic := '0';
    x_000038_000000 : std_logic := '0';
    x_000039_000000 : std_logic := '0';
    x_000040_000000 : std_logic := '0';
    x_000041_000000 : std_logic := '0';
    x_000042_000000 : std_logic := '0';
    x_000043_000000 : std_logic := '0';
    x_000044_000000 : std_logic := '0';
    x_000045_000000 : std_logic := '0';
    x_000046_000000 : std_logic := '0';
    x_000047_000000 : std_logic := '0';
    x_000048_000000 : std_logic := '0';
    x_000049_000000 : std_logic := '0';
    x_000050_000000 : std_logic := '0';
    x_000051_000000 : std_logic := '0';
    x_000052_000000 : std_logic := '0';
    x_000053_000000 : std_logic := '0';
    x_000054_000000 : std_logic := '0';
    x_000055_000000 : std_logic := '0';
    x_000056_000000 : std_logic := '0';
    x_000057_000000 : std_logic := '0';
    x_000058_000000 : std_logic := '0';
    x_000059_000000 : std_logic := '0';
    x_000060_000000 : std_logic := '0';
    x_000061_000000 : std_logic := '0';
    x_000062_000000 : std_logic := '0';
    x_000063_000000 : std_logic := '0';
    x_000064_000000 : std_logic := '0';
    x_000065_000000 : std_logic := '0';
    x_000066_000000 : std_logic := '0';
    x_000067_000000 : std_logic := '0';
    x_000068_000000 : std_logic := '0';
    x_000069_000000 : std_logic := '0';
    x_000070_000000 : std_logic := '0';
    x_000071_000000 : std_logic := '0';
    x_000072_000000 : std_logic := '0';
    x_000073_000000 : std_logic := '0';
    x_000074_000000 : std_logic := '0';
    x_000075_000000 : std_logic := '0';
    x_000076_000000 : std_logic := '0';
    x_000077_000000 : std_logic := '0';
    x_000078_000000 : std_logic := '0';
    x_000079_000000 : std_logic := '0';
    x_000080_000000 : std_logic := '0';
    x_000081_000000 : std_logic := '0';
    x_000082_000000 : std_logic := '0';
    x_000083_000000 : std_logic := '0';
    x_000084_000000 : std_logic := '0';
    x_000085_000000 : std_logic := '0';
    x_000086_000000 : std_logic := '0';
    x_000087_000000 : std_logic := '0';
    x_000088_000000 : std_logic := '0';
    x_000089_000000 : std_logic := '0';
    x_000090_000000 : std_logic := '0';
    x_000091_000000 : std_logic := '0';
    x_000092_000000 : std_logic := '0';
    x_000093_000000 : std_logic := '0';
    x_000094_000000 : std_logic := '0';
    x_000095_000000 : std_logic := '0';
    x_000096_000000 : std_logic := '0';
    x_000097_000000 : std_logic := '0';
    x_000098_000000 : std_logic := '0';
    x_000099_000000 : std_logic := '0';
    x_000100_000000 : std_logic := '0';
    x_000101_000000 : std_logic := '0';
    x_000102_000000 : std_logic := '0';
    x_000103_000000 : std_logic := '0';
    x_000104_000000 : std_logic := '0';
    x_000105_000000 : std_logic := '0';
    x_000106_000000 : std_logic := '0';
    x_000107_000000 : std_logic := '0';
    x_000108_000000 : std_logic := '0';
    x_000109_000000 : std_logic := '0';
    x_000110_000000 : std_logic := '0';
    x_000111_000000 : std_logic := '0';
    x_000112_000000 : std_logic := '0';
    x_000113_000000 : std_logic := '0';
    x_000114_000000 : std_logic := '0';
    x_000115_000000 : std_logic := '0';
    x_000116_000000 : std_logic := '0';
    x_000117_000000 : std_logic := '0';
    x_000118_000000 : std_logic := '0';
    x_000119_000000 : std_logic := '0';
    x_000120_000000 : std_logic := '0';
    x_000121_000000 : std_logic := '0';
    x_000122_000000 : std_logic := '0';
    x_000123_000000 : std_logic := '0';
    x_000124_000000 : std_logic := '0';
    x_000125_000000 : std_logic := '0';
    x_000126_000000 : std_logic := '0';
    x_000127_000000 : std_logic := '0') return std_logic;

end package SingleCyclePipelinedFunctions;


package body SingleCyclePipelinedFunctions is


function large_and (
    x_000000_000000 : std_logic;
    x_000001_000000 : std_logic := '0';
    x_000002_000000 : std_logic := '0';
    x_000003_000000 : std_logic := '0';
    x_000004_000000 : std_logic := '0';
    x_000005_000000 : std_logic := '0';
    x_000006_000000 : std_logic := '0';
    x_000007_000000 : std_logic := '0';
    x_000008_000000 : std_logic := '0';
    x_000009_000000 : std_logic := '0';
    x_000010_000000 : std_logic := '0';
    x_000011_000000 : std_logic := '0';
    x_000012_000000 : std_logic := '0';
    x_000013_000000 : std_logic := '0';
    x_000014_000000 : std_logic := '0';
    x_000015_000000 : std_logic := '0';
    x_000016_000000 : std_logic := '0';
    x_000017_000000 : std_logic := '0';
    x_000018_000000 : std_logic := '0';
    x_000019_000000 : std_logic := '0';
    x_000020_000000 : std_logic := '0';
    x_000021_000000 : std_logic := '0';
    x_000022_000000 : std_logic := '0';
    x_000023_000000 : std_logic := '0';
    x_000024_000000 : std_logic := '0';
    x_000025_000000 : std_logic := '0';
    x_000026_000000 : std_logic := '0';
    x_000027_000000 : std_logic := '0';
    x_000028_000000 : std_logic := '0';
    x_000029_000000 : std_logic := '0';
    x_000030_000000 : std_logic := '0';
    x_000031_000000 : std_logic := '0';
    x_000032_000000 : std_logic := '0';
    x_000033_000000 : std_logic := '0';
    x_000034_000000 : std_logic := '0';
    x_000035_000000 : std_logic := '0';
    x_000036_000000 : std_logic := '0';
    x_000037_000000 : std_logic := '0';
    x_000038_000000 : std_logic := '0';
    x_000039_000000 : std_logic := '0';
    x_000040_000000 : std_logic := '0';
    x_000041_000000 : std_logic := '0';
    x_000042_000000 : std_logic := '0';
    x_000043_000000 : std_logic := '0';
    x_000044_000000 : std_logic := '0';
    x_000045_000000 : std_logic := '0';
    x_000046_000000 : std_logic := '0';
    x_000047_000000 : std_logic := '0';
    x_000048_000000 : std_logic := '0';
    x_000049_000000 : std_logic := '0';
    x_000050_000000 : std_logic := '0';
    x_000051_000000 : std_logic := '0';
    x_000052_000000 : std_logic := '0';
    x_000053_000000 : std_logic := '0';
    x_000054_000000 : std_logic := '0';
    x_000055_000000 : std_logic := '0';
    x_000056_000000 : std_logic := '0';
    x_000057_000000 : std_logic := '0';
    x_000058_000000 : std_logic := '0';
    x_000059_000000 : std_logic := '0';
    x_000060_000000 : std_logic := '0';
    x_000061_000000 : std_logic := '0';
    x_000062_000000 : std_logic := '0';
    x_000063_000000 : std_logic := '0';
    x_000064_000000 : std_logic := '0';
    x_000065_000000 : std_logic := '0';
    x_000066_000000 : std_logic := '0';
    x_000067_000000 : std_logic := '0';
    x_000068_000000 : std_logic := '0';
    x_000069_000000 : std_logic := '0';
    x_000070_000000 : std_logic := '0';
    x_000071_000000 : std_logic := '0';
    x_000072_000000 : std_logic := '0';
    x_000073_000000 : std_logic := '0';
    x_000074_000000 : std_logic := '0';
    x_000075_000000 : std_logic := '0';
    x_000076_000000 : std_logic := '0';
    x_000077_000000 : std_logic := '0';
    x_000078_000000 : std_logic := '0';
    x_000079_000000 : std_logic := '0';
    x_000080_000000 : std_logic := '0';
    x_000081_000000 : std_logic := '0';
    x_000082_000000 : std_logic := '0';
    x_000083_000000 : std_logic := '0';
    x_000084_000000 : std_logic := '0';
    x_000085_000000 : std_logic := '0';
    x_000086_000000 : std_logic := '0';
    x_000087_000000 : std_logic := '0';
    x_000088_000000 : std_logic := '0';
    x_000089_000000 : std_logic := '0';
    x_000090_000000 : std_logic := '0';
    x_000091_000000 : std_logic := '0';
    x_000092_000000 : std_logic := '0';
    x_000093_000000 : std_logic := '0';
    x_000094_000000 : std_logic := '0';
    x_000095_000000 : std_logic := '0';
    x_000096_000000 : std_logic := '0';
    x_000097_000000 : std_logic := '0';
    x_000098_000000 : std_logic := '0';
    x_000099_000000 : std_logic := '0';
    x_000100_000000 : std_logic := '0';
    x_000101_000000 : std_logic := '0';
    x_000102_000000 : std_logic := '0';
    x_000103_000000 : std_logic := '0';
    x_000104_000000 : std_logic := '0';
    x_000105_000000 : std_logic := '0';
    x_000106_000000 : std_logic := '0';
    x_000107_000000 : std_logic := '0';
    x_000108_000000 : std_logic := '0';
    x_000109_000000 : std_logic := '0';
    x_000110_000000 : std_logic := '0';
    x_000111_000000 : std_logic := '0';
    x_000112_000000 : std_logic := '0';
    x_000113_000000 : std_logic := '0';
    x_000114_000000 : std_logic := '0';
    x_000115_000000 : std_logic := '0';
    x_000116_000000 : std_logic := '0';
    x_000117_000000 : std_logic := '0';
    x_000118_000000 : std_logic := '0';
    x_000119_000000 : std_logic := '0';
    x_000120_000000 : std_logic := '0';
    x_000121_000000 : std_logic := '0';
    x_000122_000000 : std_logic := '0';
    x_000123_000000 : std_logic := '0';
    x_000124_000000 : std_logic := '0';
    x_000125_000000 : std_logic := '0';
    x_000126_000000 : std_logic := '0';
    x_000127_000000 : std_logic := '0') return std_logic is 

    variable x_000000_000001 : std_logic;
    variable x_000001_000001 : std_logic;
    variable x_000002_000001 : std_logic;
    variable x_000003_000001 : std_logic;
    variable x_000004_000001 : std_logic;
    variable x_000005_000001 : std_logic;
    variable x_000006_000001 : std_logic;
    variable x_000007_000001 : std_logic;
    variable x_000008_000001 : std_logic;
    variable x_000009_000001 : std_logic;
    variable x_000010_000001 : std_logic;
    variable x_000011_000001 : std_logic;
    variable x_000012_000001 : std_logic;
    variable x_000013_000001 : std_logic;
    variable x_000014_000001 : std_logic;
    variable x_000015_000001 : std_logic;
    variable x_000016_000001 : std_logic;
    variable x_000017_000001 : std_logic;
    variable x_000018_000001 : std_logic;
    variable x_000019_000001 : std_logic;
    variable x_000020_000001 : std_logic;
    variable x_000021_000001 : std_logic;
    variable x_000022_000001 : std_logic;
    variable x_000023_000001 : std_logic;
    variable x_000024_000001 : std_logic;
    variable x_000025_000001 : std_logic;
    variable x_000000_000002 : std_logic;
    variable x_000001_000002 : std_logic;
    variable x_000002_000002 : std_logic;
    variable x_000003_000002 : std_logic;
    variable x_000004_000002 : std_logic;
    variable x_000005_000002 : std_logic;
    variable x_000000_000003 : std_logic;
    variable x_000001_000003 : std_logic;

begin 
    x_000000_000001 := and_function(x_000000_000000, x_000001_000000, x_000002_000000, x_000003_000000, x_000004_000000);
    x_000001_000001 := and_function(x_000005_000000, x_000006_000000, x_000007_000000, x_000008_000000, x_000009_000000);
    x_000002_000001 := and_function(x_000010_000000, x_000011_000000, x_000012_000000, x_000013_000000, x_000014_000000);
    x_000003_000001 := and_function(x_000015_000000, x_000016_000000, x_000017_000000, x_000018_000000, x_000019_000000);
    x_000004_000001 := and_function(x_000020_000000, x_000021_000000, x_000022_000000, x_000023_000000, x_000024_000000);
    x_000005_000001 := and_function(x_000025_000000, x_000026_000000, x_000027_000000, x_000028_000000, x_000029_000000);
    x_000006_000001 := and_function(x_000030_000000, x_000031_000000, x_000032_000000, x_000033_000000, x_000034_000000);
    x_000007_000001 := and_function(x_000035_000000, x_000036_000000, x_000037_000000, x_000038_000000, x_000039_000000);
    x_000008_000001 := and_function(x_000040_000000, x_000041_000000, x_000042_000000, x_000043_000000, x_000044_000000);
    x_000009_000001 := and_function(x_000045_000000, x_000046_000000, x_000047_000000, x_000048_000000, x_000049_000000);
    x_000010_000001 := and_function(x_000050_000000, x_000051_000000, x_000052_000000, x_000053_000000, x_000054_000000);
    x_000011_000001 := and_function(x_000055_000000, x_000056_000000, x_000057_000000, x_000058_000000, x_000059_000000);
    x_000012_000001 := and_function(x_000060_000000, x_000061_000000, x_000062_000000, x_000063_000000, x_000064_000000);
    x_000013_000001 := and_function(x_000065_000000, x_000066_000000, x_000067_000000, x_000068_000000, x_000069_000000);
    x_000014_000001 := and_function(x_000070_000000, x_000071_000000, x_000072_000000, x_000073_000000, x_000074_000000);
    x_000015_000001 := and_function(x_000075_000000, x_000076_000000, x_000077_000000, x_000078_000000, x_000079_000000);
    x_000016_000001 := and_function(x_000080_000000, x_000081_000000, x_000082_000000, x_000083_000000, x_000084_000000);
    x_000017_000001 := and_function(x_000085_000000, x_000086_000000, x_000087_000000, x_000088_000000, x_000089_000000);
    x_000018_000001 := and_function(x_000090_000000, x_000091_000000, x_000092_000000, x_000093_000000, x_000094_000000);
    x_000019_000001 := and_function(x_000095_000000, x_000096_000000, x_000097_000000, x_000098_000000, x_000099_000000);
    x_000020_000001 := and_function(x_000100_000000, x_000101_000000, x_000102_000000, x_000103_000000, x_000104_000000);
    x_000021_000001 := and_function(x_000105_000000, x_000106_000000, x_000107_000000, x_000108_000000, x_000109_000000);
    x_000022_000001 := and_function(x_000110_000000, x_000111_000000, x_000112_000000, x_000113_000000, x_000114_000000);
    x_000023_000001 := and_function(x_000115_000000, x_000116_000000, x_000117_000000, x_000118_000000, x_000119_000000);
    x_000024_000001 := and_function(x_000120_000000, x_000121_000000, x_000122_000000, x_000123_000000, x_000124_000000);
    x_000025_000001 := and_function(x_000125_000000, x_000126_000000, x_000127_000000);
    x_000000_000002 := and_function(x_000000_000001, x_000001_000001, x_000002_000001, x_000003_000001, x_000004_000001);
    x_000001_000002 := and_function(x_000005_000001, x_000006_000001, x_000007_000001, x_000008_000001, x_000009_000001);
    x_000002_000002 := and_function(x_000010_000001, x_000011_000001, x_000012_000001, x_000013_000001, x_000014_000001);
    x_000003_000002 := and_function(x_000015_000001, x_000016_000001, x_000017_000001, x_000018_000001, x_000019_000001);
    x_000004_000002 := and_function(x_000020_000001, x_000021_000001, x_000022_000001, x_000023_000001, x_000024_000001);
    x_000005_000002 := and_function(x_000025_000001);
    x_000000_000003 := and_function(x_000000_000002, x_000001_000002, x_000002_000002, x_000003_000002, x_000004_000002);
    x_000001_000003 := and_function(x_000005_000002);
    return and_function(x_000000_000003, x_000001_000003);
end function;


function large_or (
    x_000000_000000 : std_logic;
    x_000001_000000 : std_logic := '0';
    x_000002_000000 : std_logic := '0';
    x_000003_000000 : std_logic := '0';
    x_000004_000000 : std_logic := '0';
    x_000005_000000 : std_logic := '0';
    x_000006_000000 : std_logic := '0';
    x_000007_000000 : std_logic := '0';
    x_000008_000000 : std_logic := '0';
    x_000009_000000 : std_logic := '0';
    x_000010_000000 : std_logic := '0';
    x_000011_000000 : std_logic := '0';
    x_000012_000000 : std_logic := '0';
    x_000013_000000 : std_logic := '0';
    x_000014_000000 : std_logic := '0';
    x_000015_000000 : std_logic := '0';
    x_000016_000000 : std_logic := '0';
    x_000017_000000 : std_logic := '0';
    x_000018_000000 : std_logic := '0';
    x_000019_000000 : std_logic := '0';
    x_000020_000000 : std_logic := '0';
    x_000021_000000 : std_logic := '0';
    x_000022_000000 : std_logic := '0';
    x_000023_000000 : std_logic := '0';
    x_000024_000000 : std_logic := '0';
    x_000025_000000 : std_logic := '0';
    x_000026_000000 : std_logic := '0';
    x_000027_000000 : std_logic := '0';
    x_000028_000000 : std_logic := '0';
    x_000029_000000 : std_logic := '0';
    x_000030_000000 : std_logic := '0';
    x_000031_000000 : std_logic := '0';
    x_000032_000000 : std_logic := '0';
    x_000033_000000 : std_logic := '0';
    x_000034_000000 : std_logic := '0';
    x_000035_000000 : std_logic := '0';
    x_000036_000000 : std_logic := '0';
    x_000037_000000 : std_logic := '0';
    x_000038_000000 : std_logic := '0';
    x_000039_000000 : std_logic := '0';
    x_000040_000000 : std_logic := '0';
    x_000041_000000 : std_logic := '0';
    x_000042_000000 : std_logic := '0';
    x_000043_000000 : std_logic := '0';
    x_000044_000000 : std_logic := '0';
    x_000045_000000 : std_logic := '0';
    x_000046_000000 : std_logic := '0';
    x_000047_000000 : std_logic := '0';
    x_000048_000000 : std_logic := '0';
    x_000049_000000 : std_logic := '0';
    x_000050_000000 : std_logic := '0';
    x_000051_000000 : std_logic := '0';
    x_000052_000000 : std_logic := '0';
    x_000053_000000 : std_logic := '0';
    x_000054_000000 : std_logic := '0';
    x_000055_000000 : std_logic := '0';
    x_000056_000000 : std_logic := '0';
    x_000057_000000 : std_logic := '0';
    x_000058_000000 : std_logic := '0';
    x_000059_000000 : std_logic := '0';
    x_000060_000000 : std_logic := '0';
    x_000061_000000 : std_logic := '0';
    x_000062_000000 : std_logic := '0';
    x_000063_000000 : std_logic := '0';
    x_000064_000000 : std_logic := '0';
    x_000065_000000 : std_logic := '0';
    x_000066_000000 : std_logic := '0';
    x_000067_000000 : std_logic := '0';
    x_000068_000000 : std_logic := '0';
    x_000069_000000 : std_logic := '0';
    x_000070_000000 : std_logic := '0';
    x_000071_000000 : std_logic := '0';
    x_000072_000000 : std_logic := '0';
    x_000073_000000 : std_logic := '0';
    x_000074_000000 : std_logic := '0';
    x_000075_000000 : std_logic := '0';
    x_000076_000000 : std_logic := '0';
    x_000077_000000 : std_logic := '0';
    x_000078_000000 : std_logic := '0';
    x_000079_000000 : std_logic := '0';
    x_000080_000000 : std_logic := '0';
    x_000081_000000 : std_logic := '0';
    x_000082_000000 : std_logic := '0';
    x_000083_000000 : std_logic := '0';
    x_000084_000000 : std_logic := '0';
    x_000085_000000 : std_logic := '0';
    x_000086_000000 : std_logic := '0';
    x_000087_000000 : std_logic := '0';
    x_000088_000000 : std_logic := '0';
    x_000089_000000 : std_logic := '0';
    x_000090_000000 : std_logic := '0';
    x_000091_000000 : std_logic := '0';
    x_000092_000000 : std_logic := '0';
    x_000093_000000 : std_logic := '0';
    x_000094_000000 : std_logic := '0';
    x_000095_000000 : std_logic := '0';
    x_000096_000000 : std_logic := '0';
    x_000097_000000 : std_logic := '0';
    x_000098_000000 : std_logic := '0';
    x_000099_000000 : std_logic := '0';
    x_000100_000000 : std_logic := '0';
    x_000101_000000 : std_logic := '0';
    x_000102_000000 : std_logic := '0';
    x_000103_000000 : std_logic := '0';
    x_000104_000000 : std_logic := '0';
    x_000105_000000 : std_logic := '0';
    x_000106_000000 : std_logic := '0';
    x_000107_000000 : std_logic := '0';
    x_000108_000000 : std_logic := '0';
    x_000109_000000 : std_logic := '0';
    x_000110_000000 : std_logic := '0';
    x_000111_000000 : std_logic := '0';
    x_000112_000000 : std_logic := '0';
    x_000113_000000 : std_logic := '0';
    x_000114_000000 : std_logic := '0';
    x_000115_000000 : std_logic := '0';
    x_000116_000000 : std_logic := '0';
    x_000117_000000 : std_logic := '0';
    x_000118_000000 : std_logic := '0';
    x_000119_000000 : std_logic := '0';
    x_000120_000000 : std_logic := '0';
    x_000121_000000 : std_logic := '0';
    x_000122_000000 : std_logic := '0';
    x_000123_000000 : std_logic := '0';
    x_000124_000000 : std_logic := '0';
    x_000125_000000 : std_logic := '0';
    x_000126_000000 : std_logic := '0';
    x_000127_000000 : std_logic := '0') return std_logic is 

    variable x_000000_000001 : std_logic;
    variable x_000001_000001 : std_logic;
    variable x_000002_000001 : std_logic;
    variable x_000003_000001 : std_logic;
    variable x_000004_000001 : std_logic;
    variable x_000005_000001 : std_logic;
    variable x_000006_000001 : std_logic;
    variable x_000007_000001 : std_logic;
    variable x_000008_000001 : std_logic;
    variable x_000009_000001 : std_logic;
    variable x_000010_000001 : std_logic;
    variable x_000011_000001 : std_logic;
    variable x_000012_000001 : std_logic;
    variable x_000013_000001 : std_logic;
    variable x_000014_000001 : std_logic;
    variable x_000015_000001 : std_logic;
    variable x_000016_000001 : std_logic;
    variable x_000017_000001 : std_logic;
    variable x_000018_000001 : std_logic;
    variable x_000019_000001 : std_logic;
    variable x_000020_000001 : std_logic;
    variable x_000021_000001 : std_logic;
    variable x_000022_000001 : std_logic;
    variable x_000023_000001 : std_logic;
    variable x_000024_000001 : std_logic;
    variable x_000025_000001 : std_logic;
    variable x_000000_000002 : std_logic;
    variable x_000001_000002 : std_logic;
    variable x_000002_000002 : std_logic;
    variable x_000003_000002 : std_logic;
    variable x_000004_000002 : std_logic;
    variable x_000005_000002 : std_logic;
    variable x_000000_000003 : std_logic;
    variable x_000001_000003 : std_logic;

begin 
    x_000000_000001 := or_function(x_000000_000000, x_000001_000000, x_000002_000000, x_000003_000000, x_000004_000000);
    x_000001_000001 := or_function(x_000005_000000, x_000006_000000, x_000007_000000, x_000008_000000, x_000009_000000);
    x_000002_000001 := or_function(x_000010_000000, x_000011_000000, x_000012_000000, x_000013_000000, x_000014_000000);
    x_000003_000001 := or_function(x_000015_000000, x_000016_000000, x_000017_000000, x_000018_000000, x_000019_000000);
    x_000004_000001 := or_function(x_000020_000000, x_000021_000000, x_000022_000000, x_000023_000000, x_000024_000000);
    x_000005_000001 := or_function(x_000025_000000, x_000026_000000, x_000027_000000, x_000028_000000, x_000029_000000);
    x_000006_000001 := or_function(x_000030_000000, x_000031_000000, x_000032_000000, x_000033_000000, x_000034_000000);
    x_000007_000001 := or_function(x_000035_000000, x_000036_000000, x_000037_000000, x_000038_000000, x_000039_000000);
    x_000008_000001 := or_function(x_000040_000000, x_000041_000000, x_000042_000000, x_000043_000000, x_000044_000000);
    x_000009_000001 := or_function(x_000045_000000, x_000046_000000, x_000047_000000, x_000048_000000, x_000049_000000);
    x_000010_000001 := or_function(x_000050_000000, x_000051_000000, x_000052_000000, x_000053_000000, x_000054_000000);
    x_000011_000001 := or_function(x_000055_000000, x_000056_000000, x_000057_000000, x_000058_000000, x_000059_000000);
    x_000012_000001 := or_function(x_000060_000000, x_000061_000000, x_000062_000000, x_000063_000000, x_000064_000000);
    x_000013_000001 := or_function(x_000065_000000, x_000066_000000, x_000067_000000, x_000068_000000, x_000069_000000);
    x_000014_000001 := or_function(x_000070_000000, x_000071_000000, x_000072_000000, x_000073_000000, x_000074_000000);
    x_000015_000001 := or_function(x_000075_000000, x_000076_000000, x_000077_000000, x_000078_000000, x_000079_000000);
    x_000016_000001 := or_function(x_000080_000000, x_000081_000000, x_000082_000000, x_000083_000000, x_000084_000000);
    x_000017_000001 := or_function(x_000085_000000, x_000086_000000, x_000087_000000, x_000088_000000, x_000089_000000);
    x_000018_000001 := or_function(x_000090_000000, x_000091_000000, x_000092_000000, x_000093_000000, x_000094_000000);
    x_000019_000001 := or_function(x_000095_000000, x_000096_000000, x_000097_000000, x_000098_000000, x_000099_000000);
    x_000020_000001 := or_function(x_000100_000000, x_000101_000000, x_000102_000000, x_000103_000000, x_000104_000000);
    x_000021_000001 := or_function(x_000105_000000, x_000106_000000, x_000107_000000, x_000108_000000, x_000109_000000);
    x_000022_000001 := or_function(x_000110_000000, x_000111_000000, x_000112_000000, x_000113_000000, x_000114_000000);
    x_000023_000001 := or_function(x_000115_000000, x_000116_000000, x_000117_000000, x_000118_000000, x_000119_000000);
    x_000024_000001 := or_function(x_000120_000000, x_000121_000000, x_000122_000000, x_000123_000000, x_000124_000000);
    x_000025_000001 := or_function(x_000125_000000, x_000126_000000, x_000127_000000);
    x_000000_000002 := or_function(x_000000_000001, x_000001_000001, x_000002_000001, x_000003_000001, x_000004_000001);
    x_000001_000002 := or_function(x_000005_000001, x_000006_000001, x_000007_000001, x_000008_000001, x_000009_000001);
    x_000002_000002 := or_function(x_000010_000001, x_000011_000001, x_000012_000001, x_000013_000001, x_000014_000001);
    x_000003_000002 := or_function(x_000015_000001, x_000016_000001, x_000017_000001, x_000018_000001, x_000019_000001);
    x_000004_000002 := or_function(x_000020_000001, x_000021_000001, x_000022_000001, x_000023_000001, x_000024_000001);
    x_000005_000002 := or_function(x_000025_000001);
    x_000000_000003 := or_function(x_000000_000002, x_000001_000002, x_000002_000002, x_000003_000002, x_000004_000002);
    x_000001_000003 := or_function(x_000005_000002);
    return or_function(x_000000_000003, x_000001_000003);
end function;


function large_nand (
    x_000000_000000 : std_logic;
    x_000001_000000 : std_logic := '0';
    x_000002_000000 : std_logic := '0';
    x_000003_000000 : std_logic := '0';
    x_000004_000000 : std_logic := '0';
    x_000005_000000 : std_logic := '0';
    x_000006_000000 : std_logic := '0';
    x_000007_000000 : std_logic := '0';
    x_000008_000000 : std_logic := '0';
    x_000009_000000 : std_logic := '0';
    x_000010_000000 : std_logic := '0';
    x_000011_000000 : std_logic := '0';
    x_000012_000000 : std_logic := '0';
    x_000013_000000 : std_logic := '0';
    x_000014_000000 : std_logic := '0';
    x_000015_000000 : std_logic := '0';
    x_000016_000000 : std_logic := '0';
    x_000017_000000 : std_logic := '0';
    x_000018_000000 : std_logic := '0';
    x_000019_000000 : std_logic := '0';
    x_000020_000000 : std_logic := '0';
    x_000021_000000 : std_logic := '0';
    x_000022_000000 : std_logic := '0';
    x_000023_000000 : std_logic := '0';
    x_000024_000000 : std_logic := '0';
    x_000025_000000 : std_logic := '0';
    x_000026_000000 : std_logic := '0';
    x_000027_000000 : std_logic := '0';
    x_000028_000000 : std_logic := '0';
    x_000029_000000 : std_logic := '0';
    x_000030_000000 : std_logic := '0';
    x_000031_000000 : std_logic := '0';
    x_000032_000000 : std_logic := '0';
    x_000033_000000 : std_logic := '0';
    x_000034_000000 : std_logic := '0';
    x_000035_000000 : std_logic := '0';
    x_000036_000000 : std_logic := '0';
    x_000037_000000 : std_logic := '0';
    x_000038_000000 : std_logic := '0';
    x_000039_000000 : std_logic := '0';
    x_000040_000000 : std_logic := '0';
    x_000041_000000 : std_logic := '0';
    x_000042_000000 : std_logic := '0';
    x_000043_000000 : std_logic := '0';
    x_000044_000000 : std_logic := '0';
    x_000045_000000 : std_logic := '0';
    x_000046_000000 : std_logic := '0';
    x_000047_000000 : std_logic := '0';
    x_000048_000000 : std_logic := '0';
    x_000049_000000 : std_logic := '0';
    x_000050_000000 : std_logic := '0';
    x_000051_000000 : std_logic := '0';
    x_000052_000000 : std_logic := '0';
    x_000053_000000 : std_logic := '0';
    x_000054_000000 : std_logic := '0';
    x_000055_000000 : std_logic := '0';
    x_000056_000000 : std_logic := '0';
    x_000057_000000 : std_logic := '0';
    x_000058_000000 : std_logic := '0';
    x_000059_000000 : std_logic := '0';
    x_000060_000000 : std_logic := '0';
    x_000061_000000 : std_logic := '0';
    x_000062_000000 : std_logic := '0';
    x_000063_000000 : std_logic := '0';
    x_000064_000000 : std_logic := '0';
    x_000065_000000 : std_logic := '0';
    x_000066_000000 : std_logic := '0';
    x_000067_000000 : std_logic := '0';
    x_000068_000000 : std_logic := '0';
    x_000069_000000 : std_logic := '0';
    x_000070_000000 : std_logic := '0';
    x_000071_000000 : std_logic := '0';
    x_000072_000000 : std_logic := '0';
    x_000073_000000 : std_logic := '0';
    x_000074_000000 : std_logic := '0';
    x_000075_000000 : std_logic := '0';
    x_000076_000000 : std_logic := '0';
    x_000077_000000 : std_logic := '0';
    x_000078_000000 : std_logic := '0';
    x_000079_000000 : std_logic := '0';
    x_000080_000000 : std_logic := '0';
    x_000081_000000 : std_logic := '0';
    x_000082_000000 : std_logic := '0';
    x_000083_000000 : std_logic := '0';
    x_000084_000000 : std_logic := '0';
    x_000085_000000 : std_logic := '0';
    x_000086_000000 : std_logic := '0';
    x_000087_000000 : std_logic := '0';
    x_000088_000000 : std_logic := '0';
    x_000089_000000 : std_logic := '0';
    x_000090_000000 : std_logic := '0';
    x_000091_000000 : std_logic := '0';
    x_000092_000000 : std_logic := '0';
    x_000093_000000 : std_logic := '0';
    x_000094_000000 : std_logic := '0';
    x_000095_000000 : std_logic := '0';
    x_000096_000000 : std_logic := '0';
    x_000097_000000 : std_logic := '0';
    x_000098_000000 : std_logic := '0';
    x_000099_000000 : std_logic := '0';
    x_000100_000000 : std_logic := '0';
    x_000101_000000 : std_logic := '0';
    x_000102_000000 : std_logic := '0';
    x_000103_000000 : std_logic := '0';
    x_000104_000000 : std_logic := '0';
    x_000105_000000 : std_logic := '0';
    x_000106_000000 : std_logic := '0';
    x_000107_000000 : std_logic := '0';
    x_000108_000000 : std_logic := '0';
    x_000109_000000 : std_logic := '0';
    x_000110_000000 : std_logic := '0';
    x_000111_000000 : std_logic := '0';
    x_000112_000000 : std_logic := '0';
    x_000113_000000 : std_logic := '0';
    x_000114_000000 : std_logic := '0';
    x_000115_000000 : std_logic := '0';
    x_000116_000000 : std_logic := '0';
    x_000117_000000 : std_logic := '0';
    x_000118_000000 : std_logic := '0';
    x_000119_000000 : std_logic := '0';
    x_000120_000000 : std_logic := '0';
    x_000121_000000 : std_logic := '0';
    x_000122_000000 : std_logic := '0';
    x_000123_000000 : std_logic := '0';
    x_000124_000000 : std_logic := '0';
    x_000125_000000 : std_logic := '0';
    x_000126_000000 : std_logic := '0';
    x_000127_000000 : std_logic := '0') return std_logic is 

    variable x_000000_000001 : std_logic;
    variable x_000001_000001 : std_logic;
    variable x_000002_000001 : std_logic;
    variable x_000003_000001 : std_logic;
    variable x_000004_000001 : std_logic;
    variable x_000005_000001 : std_logic;
    variable x_000006_000001 : std_logic;
    variable x_000007_000001 : std_logic;
    variable x_000008_000001 : std_logic;
    variable x_000009_000001 : std_logic;
    variable x_000010_000001 : std_logic;
    variable x_000011_000001 : std_logic;
    variable x_000012_000001 : std_logic;
    variable x_000013_000001 : std_logic;
    variable x_000014_000001 : std_logic;
    variable x_000015_000001 : std_logic;
    variable x_000016_000001 : std_logic;
    variable x_000017_000001 : std_logic;
    variable x_000018_000001 : std_logic;
    variable x_000019_000001 : std_logic;
    variable x_000020_000001 : std_logic;
    variable x_000021_000001 : std_logic;
    variable x_000022_000001 : std_logic;
    variable x_000023_000001 : std_logic;
    variable x_000024_000001 : std_logic;
    variable x_000025_000001 : std_logic;
    variable x_000000_000002 : std_logic;
    variable x_000001_000002 : std_logic;
    variable x_000002_000002 : std_logic;
    variable x_000003_000002 : std_logic;
    variable x_000004_000002 : std_logic;
    variable x_000005_000002 : std_logic;
    variable x_000000_000003 : std_logic;
    variable x_000001_000003 : std_logic;

begin 
    x_000000_000001 := nand_function(x_000000_000000, x_000001_000000, x_000002_000000, x_000003_000000, x_000004_000000);
    x_000001_000001 := nand_function(x_000005_000000, x_000006_000000, x_000007_000000, x_000008_000000, x_000009_000000);
    x_000002_000001 := nand_function(x_000010_000000, x_000011_000000, x_000012_000000, x_000013_000000, x_000014_000000);
    x_000003_000001 := nand_function(x_000015_000000, x_000016_000000, x_000017_000000, x_000018_000000, x_000019_000000);
    x_000004_000001 := nand_function(x_000020_000000, x_000021_000000, x_000022_000000, x_000023_000000, x_000024_000000);
    x_000005_000001 := nand_function(x_000025_000000, x_000026_000000, x_000027_000000, x_000028_000000, x_000029_000000);
    x_000006_000001 := nand_function(x_000030_000000, x_000031_000000, x_000032_000000, x_000033_000000, x_000034_000000);
    x_000007_000001 := nand_function(x_000035_000000, x_000036_000000, x_000037_000000, x_000038_000000, x_000039_000000);
    x_000008_000001 := nand_function(x_000040_000000, x_000041_000000, x_000042_000000, x_000043_000000, x_000044_000000);
    x_000009_000001 := nand_function(x_000045_000000, x_000046_000000, x_000047_000000, x_000048_000000, x_000049_000000);
    x_000010_000001 := nand_function(x_000050_000000, x_000051_000000, x_000052_000000, x_000053_000000, x_000054_000000);
    x_000011_000001 := nand_function(x_000055_000000, x_000056_000000, x_000057_000000, x_000058_000000, x_000059_000000);
    x_000012_000001 := nand_function(x_000060_000000, x_000061_000000, x_000062_000000, x_000063_000000, x_000064_000000);
    x_000013_000001 := nand_function(x_000065_000000, x_000066_000000, x_000067_000000, x_000068_000000, x_000069_000000);
    x_000014_000001 := nand_function(x_000070_000000, x_000071_000000, x_000072_000000, x_000073_000000, x_000074_000000);
    x_000015_000001 := nand_function(x_000075_000000, x_000076_000000, x_000077_000000, x_000078_000000, x_000079_000000);
    x_000016_000001 := nand_function(x_000080_000000, x_000081_000000, x_000082_000000, x_000083_000000, x_000084_000000);
    x_000017_000001 := nand_function(x_000085_000000, x_000086_000000, x_000087_000000, x_000088_000000, x_000089_000000);
    x_000018_000001 := nand_function(x_000090_000000, x_000091_000000, x_000092_000000, x_000093_000000, x_000094_000000);
    x_000019_000001 := nand_function(x_000095_000000, x_000096_000000, x_000097_000000, x_000098_000000, x_000099_000000);
    x_000020_000001 := nand_function(x_000100_000000, x_000101_000000, x_000102_000000, x_000103_000000, x_000104_000000);
    x_000021_000001 := nand_function(x_000105_000000, x_000106_000000, x_000107_000000, x_000108_000000, x_000109_000000);
    x_000022_000001 := nand_function(x_000110_000000, x_000111_000000, x_000112_000000, x_000113_000000, x_000114_000000);
    x_000023_000001 := nand_function(x_000115_000000, x_000116_000000, x_000117_000000, x_000118_000000, x_000119_000000);
    x_000024_000001 := nand_function(x_000120_000000, x_000121_000000, x_000122_000000, x_000123_000000, x_000124_000000);
    x_000025_000001 := nand_function(x_000125_000000, x_000126_000000, x_000127_000000);
    x_000000_000002 := nand_function(x_000000_000001, x_000001_000001, x_000002_000001, x_000003_000001, x_000004_000001);
    x_000001_000002 := nand_function(x_000005_000001, x_000006_000001, x_000007_000001, x_000008_000001, x_000009_000001);
    x_000002_000002 := nand_function(x_000010_000001, x_000011_000001, x_000012_000001, x_000013_000001, x_000014_000001);
    x_000003_000002 := nand_function(x_000015_000001, x_000016_000001, x_000017_000001, x_000018_000001, x_000019_000001);
    x_000004_000002 := nand_function(x_000020_000001, x_000021_000001, x_000022_000001, x_000023_000001, x_000024_000001);
    x_000005_000002 := nand_function(x_000025_000001);
    x_000000_000003 := nand_function(x_000000_000002, x_000001_000002, x_000002_000002, x_000003_000002, x_000004_000002);
    x_000001_000003 := nand_function(x_000005_000002);
    return nand_function(x_000000_000003, x_000001_000003);
end function;


function large_nor (
    x_000000_000000 : std_logic;
    x_000001_000000 : std_logic := '0';
    x_000002_000000 : std_logic := '0';
    x_000003_000000 : std_logic := '0';
    x_000004_000000 : std_logic := '0';
    x_000005_000000 : std_logic := '0';
    x_000006_000000 : std_logic := '0';
    x_000007_000000 : std_logic := '0';
    x_000008_000000 : std_logic := '0';
    x_000009_000000 : std_logic := '0';
    x_000010_000000 : std_logic := '0';
    x_000011_000000 : std_logic := '0';
    x_000012_000000 : std_logic := '0';
    x_000013_000000 : std_logic := '0';
    x_000014_000000 : std_logic := '0';
    x_000015_000000 : std_logic := '0';
    x_000016_000000 : std_logic := '0';
    x_000017_000000 : std_logic := '0';
    x_000018_000000 : std_logic := '0';
    x_000019_000000 : std_logic := '0';
    x_000020_000000 : std_logic := '0';
    x_000021_000000 : std_logic := '0';
    x_000022_000000 : std_logic := '0';
    x_000023_000000 : std_logic := '0';
    x_000024_000000 : std_logic := '0';
    x_000025_000000 : std_logic := '0';
    x_000026_000000 : std_logic := '0';
    x_000027_000000 : std_logic := '0';
    x_000028_000000 : std_logic := '0';
    x_000029_000000 : std_logic := '0';
    x_000030_000000 : std_logic := '0';
    x_000031_000000 : std_logic := '0';
    x_000032_000000 : std_logic := '0';
    x_000033_000000 : std_logic := '0';
    x_000034_000000 : std_logic := '0';
    x_000035_000000 : std_logic := '0';
    x_000036_000000 : std_logic := '0';
    x_000037_000000 : std_logic := '0';
    x_000038_000000 : std_logic := '0';
    x_000039_000000 : std_logic := '0';
    x_000040_000000 : std_logic := '0';
    x_000041_000000 : std_logic := '0';
    x_000042_000000 : std_logic := '0';
    x_000043_000000 : std_logic := '0';
    x_000044_000000 : std_logic := '0';
    x_000045_000000 : std_logic := '0';
    x_000046_000000 : std_logic := '0';
    x_000047_000000 : std_logic := '0';
    x_000048_000000 : std_logic := '0';
    x_000049_000000 : std_logic := '0';
    x_000050_000000 : std_logic := '0';
    x_000051_000000 : std_logic := '0';
    x_000052_000000 : std_logic := '0';
    x_000053_000000 : std_logic := '0';
    x_000054_000000 : std_logic := '0';
    x_000055_000000 : std_logic := '0';
    x_000056_000000 : std_logic := '0';
    x_000057_000000 : std_logic := '0';
    x_000058_000000 : std_logic := '0';
    x_000059_000000 : std_logic := '0';
    x_000060_000000 : std_logic := '0';
    x_000061_000000 : std_logic := '0';
    x_000062_000000 : std_logic := '0';
    x_000063_000000 : std_logic := '0';
    x_000064_000000 : std_logic := '0';
    x_000065_000000 : std_logic := '0';
    x_000066_000000 : std_logic := '0';
    x_000067_000000 : std_logic := '0';
    x_000068_000000 : std_logic := '0';
    x_000069_000000 : std_logic := '0';
    x_000070_000000 : std_logic := '0';
    x_000071_000000 : std_logic := '0';
    x_000072_000000 : std_logic := '0';
    x_000073_000000 : std_logic := '0';
    x_000074_000000 : std_logic := '0';
    x_000075_000000 : std_logic := '0';
    x_000076_000000 : std_logic := '0';
    x_000077_000000 : std_logic := '0';
    x_000078_000000 : std_logic := '0';
    x_000079_000000 : std_logic := '0';
    x_000080_000000 : std_logic := '0';
    x_000081_000000 : std_logic := '0';
    x_000082_000000 : std_logic := '0';
    x_000083_000000 : std_logic := '0';
    x_000084_000000 : std_logic := '0';
    x_000085_000000 : std_logic := '0';
    x_000086_000000 : std_logic := '0';
    x_000087_000000 : std_logic := '0';
    x_000088_000000 : std_logic := '0';
    x_000089_000000 : std_logic := '0';
    x_000090_000000 : std_logic := '0';
    x_000091_000000 : std_logic := '0';
    x_000092_000000 : std_logic := '0';
    x_000093_000000 : std_logic := '0';
    x_000094_000000 : std_logic := '0';
    x_000095_000000 : std_logic := '0';
    x_000096_000000 : std_logic := '0';
    x_000097_000000 : std_logic := '0';
    x_000098_000000 : std_logic := '0';
    x_000099_000000 : std_logic := '0';
    x_000100_000000 : std_logic := '0';
    x_000101_000000 : std_logic := '0';
    x_000102_000000 : std_logic := '0';
    x_000103_000000 : std_logic := '0';
    x_000104_000000 : std_logic := '0';
    x_000105_000000 : std_logic := '0';
    x_000106_000000 : std_logic := '0';
    x_000107_000000 : std_logic := '0';
    x_000108_000000 : std_logic := '0';
    x_000109_000000 : std_logic := '0';
    x_000110_000000 : std_logic := '0';
    x_000111_000000 : std_logic := '0';
    x_000112_000000 : std_logic := '0';
    x_000113_000000 : std_logic := '0';
    x_000114_000000 : std_logic := '0';
    x_000115_000000 : std_logic := '0';
    x_000116_000000 : std_logic := '0';
    x_000117_000000 : std_logic := '0';
    x_000118_000000 : std_logic := '0';
    x_000119_000000 : std_logic := '0';
    x_000120_000000 : std_logic := '0';
    x_000121_000000 : std_logic := '0';
    x_000122_000000 : std_logic := '0';
    x_000123_000000 : std_logic := '0';
    x_000124_000000 : std_logic := '0';
    x_000125_000000 : std_logic := '0';
    x_000126_000000 : std_logic := '0';
    x_000127_000000 : std_logic := '0') return std_logic is 

    variable x_000000_000001 : std_logic;
    variable x_000001_000001 : std_logic;
    variable x_000002_000001 : std_logic;
    variable x_000003_000001 : std_logic;
    variable x_000004_000001 : std_logic;
    variable x_000005_000001 : std_logic;
    variable x_000006_000001 : std_logic;
    variable x_000007_000001 : std_logic;
    variable x_000008_000001 : std_logic;
    variable x_000009_000001 : std_logic;
    variable x_000010_000001 : std_logic;
    variable x_000011_000001 : std_logic;
    variable x_000012_000001 : std_logic;
    variable x_000013_000001 : std_logic;
    variable x_000014_000001 : std_logic;
    variable x_000015_000001 : std_logic;
    variable x_000016_000001 : std_logic;
    variable x_000017_000001 : std_logic;
    variable x_000018_000001 : std_logic;
    variable x_000019_000001 : std_logic;
    variable x_000020_000001 : std_logic;
    variable x_000021_000001 : std_logic;
    variable x_000022_000001 : std_logic;
    variable x_000023_000001 : std_logic;
    variable x_000024_000001 : std_logic;
    variable x_000025_000001 : std_logic;
    variable x_000000_000002 : std_logic;
    variable x_000001_000002 : std_logic;
    variable x_000002_000002 : std_logic;
    variable x_000003_000002 : std_logic;
    variable x_000004_000002 : std_logic;
    variable x_000005_000002 : std_logic;
    variable x_000000_000003 : std_logic;
    variable x_000001_000003 : std_logic;

begin 
    x_000000_000001 := nor_function(x_000000_000000, x_000001_000000, x_000002_000000, x_000003_000000, x_000004_000000);
    x_000001_000001 := nor_function(x_000005_000000, x_000006_000000, x_000007_000000, x_000008_000000, x_000009_000000);
    x_000002_000001 := nor_function(x_000010_000000, x_000011_000000, x_000012_000000, x_000013_000000, x_000014_000000);
    x_000003_000001 := nor_function(x_000015_000000, x_000016_000000, x_000017_000000, x_000018_000000, x_000019_000000);
    x_000004_000001 := nor_function(x_000020_000000, x_000021_000000, x_000022_000000, x_000023_000000, x_000024_000000);
    x_000005_000001 := nor_function(x_000025_000000, x_000026_000000, x_000027_000000, x_000028_000000, x_000029_000000);
    x_000006_000001 := nor_function(x_000030_000000, x_000031_000000, x_000032_000000, x_000033_000000, x_000034_000000);
    x_000007_000001 := nor_function(x_000035_000000, x_000036_000000, x_000037_000000, x_000038_000000, x_000039_000000);
    x_000008_000001 := nor_function(x_000040_000000, x_000041_000000, x_000042_000000, x_000043_000000, x_000044_000000);
    x_000009_000001 := nor_function(x_000045_000000, x_000046_000000, x_000047_000000, x_000048_000000, x_000049_000000);
    x_000010_000001 := nor_function(x_000050_000000, x_000051_000000, x_000052_000000, x_000053_000000, x_000054_000000);
    x_000011_000001 := nor_function(x_000055_000000, x_000056_000000, x_000057_000000, x_000058_000000, x_000059_000000);
    x_000012_000001 := nor_function(x_000060_000000, x_000061_000000, x_000062_000000, x_000063_000000, x_000064_000000);
    x_000013_000001 := nor_function(x_000065_000000, x_000066_000000, x_000067_000000, x_000068_000000, x_000069_000000);
    x_000014_000001 := nor_function(x_000070_000000, x_000071_000000, x_000072_000000, x_000073_000000, x_000074_000000);
    x_000015_000001 := nor_function(x_000075_000000, x_000076_000000, x_000077_000000, x_000078_000000, x_000079_000000);
    x_000016_000001 := nor_function(x_000080_000000, x_000081_000000, x_000082_000000, x_000083_000000, x_000084_000000);
    x_000017_000001 := nor_function(x_000085_000000, x_000086_000000, x_000087_000000, x_000088_000000, x_000089_000000);
    x_000018_000001 := nor_function(x_000090_000000, x_000091_000000, x_000092_000000, x_000093_000000, x_000094_000000);
    x_000019_000001 := nor_function(x_000095_000000, x_000096_000000, x_000097_000000, x_000098_000000, x_000099_000000);
    x_000020_000001 := nor_function(x_000100_000000, x_000101_000000, x_000102_000000, x_000103_000000, x_000104_000000);
    x_000021_000001 := nor_function(x_000105_000000, x_000106_000000, x_000107_000000, x_000108_000000, x_000109_000000);
    x_000022_000001 := nor_function(x_000110_000000, x_000111_000000, x_000112_000000, x_000113_000000, x_000114_000000);
    x_000023_000001 := nor_function(x_000115_000000, x_000116_000000, x_000117_000000, x_000118_000000, x_000119_000000);
    x_000024_000001 := nor_function(x_000120_000000, x_000121_000000, x_000122_000000, x_000123_000000, x_000124_000000);
    x_000025_000001 := nor_function(x_000125_000000, x_000126_000000, x_000127_000000);
    x_000000_000002 := nor_function(x_000000_000001, x_000001_000001, x_000002_000001, x_000003_000001, x_000004_000001);
    x_000001_000002 := nor_function(x_000005_000001, x_000006_000001, x_000007_000001, x_000008_000001, x_000009_000001);
    x_000002_000002 := nor_function(x_000010_000001, x_000011_000001, x_000012_000001, x_000013_000001, x_000014_000001);
    x_000003_000002 := nor_function(x_000015_000001, x_000016_000001, x_000017_000001, x_000018_000001, x_000019_000001);
    x_000004_000002 := nor_function(x_000020_000001, x_000021_000001, x_000022_000001, x_000023_000001, x_000024_000001);
    x_000005_000002 := nor_function(x_000025_000001);
    x_000000_000003 := nor_function(x_000000_000002, x_000001_000002, x_000002_000002, x_000003_000002, x_000004_000002);
    x_000001_000003 := nor_function(x_000005_000002);
    return nor_function(x_000000_000003, x_000001_000003);
end function;


function large_xor (
    x_000000_000000 : std_logic;
    x_000001_000000 : std_logic := '0';
    x_000002_000000 : std_logic := '0';
    x_000003_000000 : std_logic := '0';
    x_000004_000000 : std_logic := '0';
    x_000005_000000 : std_logic := '0';
    x_000006_000000 : std_logic := '0';
    x_000007_000000 : std_logic := '0';
    x_000008_000000 : std_logic := '0';
    x_000009_000000 : std_logic := '0';
    x_000010_000000 : std_logic := '0';
    x_000011_000000 : std_logic := '0';
    x_000012_000000 : std_logic := '0';
    x_000013_000000 : std_logic := '0';
    x_000014_000000 : std_logic := '0';
    x_000015_000000 : std_logic := '0';
    x_000016_000000 : std_logic := '0';
    x_000017_000000 : std_logic := '0';
    x_000018_000000 : std_logic := '0';
    x_000019_000000 : std_logic := '0';
    x_000020_000000 : std_logic := '0';
    x_000021_000000 : std_logic := '0';
    x_000022_000000 : std_logic := '0';
    x_000023_000000 : std_logic := '0';
    x_000024_000000 : std_logic := '0';
    x_000025_000000 : std_logic := '0';
    x_000026_000000 : std_logic := '0';
    x_000027_000000 : std_logic := '0';
    x_000028_000000 : std_logic := '0';
    x_000029_000000 : std_logic := '0';
    x_000030_000000 : std_logic := '0';
    x_000031_000000 : std_logic := '0';
    x_000032_000000 : std_logic := '0';
    x_000033_000000 : std_logic := '0';
    x_000034_000000 : std_logic := '0';
    x_000035_000000 : std_logic := '0';
    x_000036_000000 : std_logic := '0';
    x_000037_000000 : std_logic := '0';
    x_000038_000000 : std_logic := '0';
    x_000039_000000 : std_logic := '0';
    x_000040_000000 : std_logic := '0';
    x_000041_000000 : std_logic := '0';
    x_000042_000000 : std_logic := '0';
    x_000043_000000 : std_logic := '0';
    x_000044_000000 : std_logic := '0';
    x_000045_000000 : std_logic := '0';
    x_000046_000000 : std_logic := '0';
    x_000047_000000 : std_logic := '0';
    x_000048_000000 : std_logic := '0';
    x_000049_000000 : std_logic := '0';
    x_000050_000000 : std_logic := '0';
    x_000051_000000 : std_logic := '0';
    x_000052_000000 : std_logic := '0';
    x_000053_000000 : std_logic := '0';
    x_000054_000000 : std_logic := '0';
    x_000055_000000 : std_logic := '0';
    x_000056_000000 : std_logic := '0';
    x_000057_000000 : std_logic := '0';
    x_000058_000000 : std_logic := '0';
    x_000059_000000 : std_logic := '0';
    x_000060_000000 : std_logic := '0';
    x_000061_000000 : std_logic := '0';
    x_000062_000000 : std_logic := '0';
    x_000063_000000 : std_logic := '0';
    x_000064_000000 : std_logic := '0';
    x_000065_000000 : std_logic := '0';
    x_000066_000000 : std_logic := '0';
    x_000067_000000 : std_logic := '0';
    x_000068_000000 : std_logic := '0';
    x_000069_000000 : std_logic := '0';
    x_000070_000000 : std_logic := '0';
    x_000071_000000 : std_logic := '0';
    x_000072_000000 : std_logic := '0';
    x_000073_000000 : std_logic := '0';
    x_000074_000000 : std_logic := '0';
    x_000075_000000 : std_logic := '0';
    x_000076_000000 : std_logic := '0';
    x_000077_000000 : std_logic := '0';
    x_000078_000000 : std_logic := '0';
    x_000079_000000 : std_logic := '0';
    x_000080_000000 : std_logic := '0';
    x_000081_000000 : std_logic := '0';
    x_000082_000000 : std_logic := '0';
    x_000083_000000 : std_logic := '0';
    x_000084_000000 : std_logic := '0';
    x_000085_000000 : std_logic := '0';
    x_000086_000000 : std_logic := '0';
    x_000087_000000 : std_logic := '0';
    x_000088_000000 : std_logic := '0';
    x_000089_000000 : std_logic := '0';
    x_000090_000000 : std_logic := '0';
    x_000091_000000 : std_logic := '0';
    x_000092_000000 : std_logic := '0';
    x_000093_000000 : std_logic := '0';
    x_000094_000000 : std_logic := '0';
    x_000095_000000 : std_logic := '0';
    x_000096_000000 : std_logic := '0';
    x_000097_000000 : std_logic := '0';
    x_000098_000000 : std_logic := '0';
    x_000099_000000 : std_logic := '0';
    x_000100_000000 : std_logic := '0';
    x_000101_000000 : std_logic := '0';
    x_000102_000000 : std_logic := '0';
    x_000103_000000 : std_logic := '0';
    x_000104_000000 : std_logic := '0';
    x_000105_000000 : std_logic := '0';
    x_000106_000000 : std_logic := '0';
    x_000107_000000 : std_logic := '0';
    x_000108_000000 : std_logic := '0';
    x_000109_000000 : std_logic := '0';
    x_000110_000000 : std_logic := '0';
    x_000111_000000 : std_logic := '0';
    x_000112_000000 : std_logic := '0';
    x_000113_000000 : std_logic := '0';
    x_000114_000000 : std_logic := '0';
    x_000115_000000 : std_logic := '0';
    x_000116_000000 : std_logic := '0';
    x_000117_000000 : std_logic := '0';
    x_000118_000000 : std_logic := '0';
    x_000119_000000 : std_logic := '0';
    x_000120_000000 : std_logic := '0';
    x_000121_000000 : std_logic := '0';
    x_000122_000000 : std_logic := '0';
    x_000123_000000 : std_logic := '0';
    x_000124_000000 : std_logic := '0';
    x_000125_000000 : std_logic := '0';
    x_000126_000000 : std_logic := '0';
    x_000127_000000 : std_logic := '0') return std_logic is 

    variable x_000000_000001 : std_logic;
    variable x_000001_000001 : std_logic;
    variable x_000002_000001 : std_logic;
    variable x_000003_000001 : std_logic;
    variable x_000004_000001 : std_logic;
    variable x_000005_000001 : std_logic;
    variable x_000006_000001 : std_logic;
    variable x_000007_000001 : std_logic;
    variable x_000008_000001 : std_logic;
    variable x_000009_000001 : std_logic;
    variable x_000010_000001 : std_logic;
    variable x_000011_000001 : std_logic;
    variable x_000012_000001 : std_logic;
    variable x_000013_000001 : std_logic;
    variable x_000014_000001 : std_logic;
    variable x_000015_000001 : std_logic;
    variable x_000016_000001 : std_logic;
    variable x_000017_000001 : std_logic;
    variable x_000018_000001 : std_logic;
    variable x_000019_000001 : std_logic;
    variable x_000020_000001 : std_logic;
    variable x_000021_000001 : std_logic;
    variable x_000022_000001 : std_logic;
    variable x_000023_000001 : std_logic;
    variable x_000024_000001 : std_logic;
    variable x_000025_000001 : std_logic;
    variable x_000000_000002 : std_logic;
    variable x_000001_000002 : std_logic;
    variable x_000002_000002 : std_logic;
    variable x_000003_000002 : std_logic;
    variable x_000004_000002 : std_logic;
    variable x_000005_000002 : std_logic;
    variable x_000000_000003 : std_logic;
    variable x_000001_000003 : std_logic;

begin 
    x_000000_000001 := xor_function(x_000000_000000, x_000001_000000, x_000002_000000, x_000003_000000, x_000004_000000);
    x_000001_000001 := xor_function(x_000005_000000, x_000006_000000, x_000007_000000, x_000008_000000, x_000009_000000);
    x_000002_000001 := xor_function(x_000010_000000, x_000011_000000, x_000012_000000, x_000013_000000, x_000014_000000);
    x_000003_000001 := xor_function(x_000015_000000, x_000016_000000, x_000017_000000, x_000018_000000, x_000019_000000);
    x_000004_000001 := xor_function(x_000020_000000, x_000021_000000, x_000022_000000, x_000023_000000, x_000024_000000);
    x_000005_000001 := xor_function(x_000025_000000, x_000026_000000, x_000027_000000, x_000028_000000, x_000029_000000);
    x_000006_000001 := xor_function(x_000030_000000, x_000031_000000, x_000032_000000, x_000033_000000, x_000034_000000);
    x_000007_000001 := xor_function(x_000035_000000, x_000036_000000, x_000037_000000, x_000038_000000, x_000039_000000);
    x_000008_000001 := xor_function(x_000040_000000, x_000041_000000, x_000042_000000, x_000043_000000, x_000044_000000);
    x_000009_000001 := xor_function(x_000045_000000, x_000046_000000, x_000047_000000, x_000048_000000, x_000049_000000);
    x_000010_000001 := xor_function(x_000050_000000, x_000051_000000, x_000052_000000, x_000053_000000, x_000054_000000);
    x_000011_000001 := xor_function(x_000055_000000, x_000056_000000, x_000057_000000, x_000058_000000, x_000059_000000);
    x_000012_000001 := xor_function(x_000060_000000, x_000061_000000, x_000062_000000, x_000063_000000, x_000064_000000);
    x_000013_000001 := xor_function(x_000065_000000, x_000066_000000, x_000067_000000, x_000068_000000, x_000069_000000);
    x_000014_000001 := xor_function(x_000070_000000, x_000071_000000, x_000072_000000, x_000073_000000, x_000074_000000);
    x_000015_000001 := xor_function(x_000075_000000, x_000076_000000, x_000077_000000, x_000078_000000, x_000079_000000);
    x_000016_000001 := xor_function(x_000080_000000, x_000081_000000, x_000082_000000, x_000083_000000, x_000084_000000);
    x_000017_000001 := xor_function(x_000085_000000, x_000086_000000, x_000087_000000, x_000088_000000, x_000089_000000);
    x_000018_000001 := xor_function(x_000090_000000, x_000091_000000, x_000092_000000, x_000093_000000, x_000094_000000);
    x_000019_000001 := xor_function(x_000095_000000, x_000096_000000, x_000097_000000, x_000098_000000, x_000099_000000);
    x_000020_000001 := xor_function(x_000100_000000, x_000101_000000, x_000102_000000, x_000103_000000, x_000104_000000);
    x_000021_000001 := xor_function(x_000105_000000, x_000106_000000, x_000107_000000, x_000108_000000, x_000109_000000);
    x_000022_000001 := xor_function(x_000110_000000, x_000111_000000, x_000112_000000, x_000113_000000, x_000114_000000);
    x_000023_000001 := xor_function(x_000115_000000, x_000116_000000, x_000117_000000, x_000118_000000, x_000119_000000);
    x_000024_000001 := xor_function(x_000120_000000, x_000121_000000, x_000122_000000, x_000123_000000, x_000124_000000);
    x_000025_000001 := xor_function(x_000125_000000, x_000126_000000, x_000127_000000);
    x_000000_000002 := xor_function(x_000000_000001, x_000001_000001, x_000002_000001, x_000003_000001, x_000004_000001);
    x_000001_000002 := xor_function(x_000005_000001, x_000006_000001, x_000007_000001, x_000008_000001, x_000009_000001);
    x_000002_000002 := xor_function(x_000010_000001, x_000011_000001, x_000012_000001, x_000013_000001, x_000014_000001);
    x_000003_000002 := xor_function(x_000015_000001, x_000016_000001, x_000017_000001, x_000018_000001, x_000019_000001);
    x_000004_000002 := xor_function(x_000020_000001, x_000021_000001, x_000022_000001, x_000023_000001, x_000024_000001);
    x_000005_000002 := xor_function(x_000025_000001);
    x_000000_000003 := xor_function(x_000000_000002, x_000001_000002, x_000002_000002, x_000003_000002, x_000004_000002);
    x_000001_000003 := xor_function(x_000005_000002);
    return xor_function(x_000000_000003, x_000001_000003);
end function;

end package body SingleCyclePipelinedFunctions;
