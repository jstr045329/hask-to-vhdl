----------------------------------------------------------------------------------------------------
--                                   Testbench for MinFunction
----------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.VhdSimToolsPkg.all;
use work.MinFunction_0016;

entity MinFunction_0064_tb is
end MinFunction_0064_tb;


architecture behavioral_MinFunction_0064_tb of MinFunction_0064_tb is


component MinFunction_0064 is 
    generic ( 
        max_integer : integer := (2**30) - 2
    );    
    port (
        clk : in std_logic;
        rst : in std_logic;
        i_soft_rst : in std_logic;
        i_distance_0000 : in integer := max_integer;
        i_distance_0001 : in integer := max_integer;
        i_distance_0002 : in integer := max_integer;
        i_distance_0003 : in integer := max_integer;
        i_distance_0004 : in integer := max_integer;
        i_distance_0005 : in integer := max_integer;
        i_distance_0006 : in integer := max_integer;
        i_distance_0007 : in integer := max_integer;
        i_distance_0008 : in integer := max_integer;
        i_distance_0009 : in integer := max_integer;
        i_distance_0010 : in integer := max_integer;
        i_distance_0011 : in integer := max_integer;
        i_distance_0012 : in integer := max_integer;
        i_distance_0013 : in integer := max_integer;
        i_distance_0014 : in integer := max_integer;
        i_distance_0015 : in integer := max_integer;
        i_distance_0016 : in integer := max_integer;
        i_distance_0017 : in integer := max_integer;
        i_distance_0018 : in integer := max_integer;
        i_distance_0019 : in integer := max_integer;
        i_distance_0020 : in integer := max_integer;
        i_distance_0021 : in integer := max_integer;
        i_distance_0022 : in integer := max_integer;
        i_distance_0023 : in integer := max_integer;
        i_distance_0024 : in integer := max_integer;
        i_distance_0025 : in integer := max_integer;
        i_distance_0026 : in integer := max_integer;
        i_distance_0027 : in integer := max_integer;
        i_distance_0028 : in integer := max_integer;
        i_distance_0029 : in integer := max_integer;
        i_distance_0030 : in integer := max_integer;
        i_distance_0031 : in integer := max_integer;
        i_distance_0032 : in integer := max_integer;
        i_distance_0033 : in integer := max_integer;
        i_distance_0034 : in integer := max_integer;
        i_distance_0035 : in integer := max_integer;
        i_distance_0036 : in integer := max_integer;
        i_distance_0037 : in integer := max_integer;
        i_distance_0038 : in integer := max_integer;
        i_distance_0039 : in integer := max_integer;
        i_distance_0040 : in integer := max_integer;
        i_distance_0041 : in integer := max_integer;
        i_distance_0042 : in integer := max_integer;
        i_distance_0043 : in integer := max_integer;
        i_distance_0044 : in integer := max_integer;
        i_distance_0045 : in integer := max_integer;
        i_distance_0046 : in integer := max_integer;
        i_distance_0047 : in integer := max_integer;
        i_distance_0048 : in integer := max_integer;
        i_distance_0049 : in integer := max_integer;
        i_distance_0050 : in integer := max_integer;
        i_distance_0051 : in integer := max_integer;
        i_distance_0052 : in integer := max_integer;
        i_distance_0053 : in integer := max_integer;
        i_distance_0054 : in integer := max_integer;
        i_distance_0055 : in integer := max_integer;
        i_distance_0056 : in integer := max_integer;
        i_distance_0057 : in integer := max_integer;
        i_distance_0058 : in integer := max_integer;
        i_distance_0059 : in integer := max_integer;
        i_distance_0060 : in integer := max_integer;
        i_distance_0061 : in integer := max_integer;
        i_distance_0062 : in integer := max_integer;
        i_distance_0063 : in integer := max_integer;
        o_min : out integer;
        o_latency : out integer
    );
end component;


signal clk : std_logic := '1';
signal rst : std_logic := '1';
signal i_soft_rst : std_logic;
signal i_distance_0000 : integer;
signal i_distance_0001 : integer;
signal i_distance_0002 : integer;
signal i_distance_0003 : integer;
signal i_distance_0004 : integer;
signal i_distance_0005 : integer;
signal i_distance_0006 : integer;
signal i_distance_0007 : integer;
signal i_distance_0008 : integer;
signal i_distance_0009 : integer;
signal i_distance_0010 : integer;
signal i_distance_0011 : integer;
signal i_distance_0012 : integer;
signal i_distance_0013 : integer;
signal i_distance_0014 : integer;
signal i_distance_0015 : integer;
signal i_distance_0016 : integer;
signal i_distance_0017 : integer;
signal i_distance_0018 : integer;
signal i_distance_0019 : integer;
signal i_distance_0020 : integer;
signal i_distance_0021 : integer;
signal i_distance_0022 : integer;
signal i_distance_0023 : integer;
signal i_distance_0024 : integer;
signal i_distance_0025 : integer;
signal i_distance_0026 : integer;
signal i_distance_0027 : integer;
signal i_distance_0028 : integer;
signal i_distance_0029 : integer;
signal i_distance_0030 : integer;
signal i_distance_0031 : integer;
signal i_distance_0032 : integer;
signal i_distance_0033 : integer;
signal i_distance_0034 : integer;
signal i_distance_0035 : integer;
signal i_distance_0036 : integer;
signal i_distance_0037 : integer;
signal i_distance_0038 : integer;
signal i_distance_0039 : integer;
signal i_distance_0040 : integer;
signal i_distance_0041 : integer;
signal i_distance_0042 : integer;
signal i_distance_0043 : integer;
signal i_distance_0044 : integer;
signal i_distance_0045 : integer;
signal i_distance_0046 : integer;
signal i_distance_0047 : integer;
signal i_distance_0048 : integer;
signal i_distance_0049 : integer;
signal i_distance_0050 : integer;
signal i_distance_0051 : integer;
signal i_distance_0052 : integer;
signal i_distance_0053 : integer;
signal i_distance_0054 : integer;
signal i_distance_0055 : integer;
signal i_distance_0056 : integer;
signal i_distance_0057 : integer;
signal i_distance_0058 : integer;
signal i_distance_0059 : integer;
signal i_distance_0060 : integer;
signal i_distance_0061 : integer;
signal i_distance_0062 : integer;
signal i_distance_0063 : integer;
signal o_min : integer;
signal o_latency : integer;

signal correct_answer : integer;

constant clk_per : time := 10 ns;
signal sim_done : std_logic := '0';
signal test_stage : integer := 0;


begin


----------------------------------------------------------------------------------------------------
--                                          Boiler Plate
----------------------------------------------------------------------------------------------------
CLOCK_PROCESS: process
begin
    if sim_done = '1' then
        wait;
    else
        wait for clk_per/2;
        clk <= not clk;
    end if;
end process;


----------------------------------------------------------------------------------------------------
--                                          Stim Process
----------------------------------------------------------------------------------------------------
STIM_PROCESS: process
begin
    i_soft_rst <= '0';
    i_distance_0000 <= (2**30)-1;
    i_distance_0001 <= (2**30)-1;
    i_distance_0002 <= (2**30)-1;
    i_distance_0003 <= (2**30)-1;
    i_distance_0004 <= (2**30)-1;
    i_distance_0005 <= (2**30)-1;
    i_distance_0006 <= (2**30)-1;
    i_distance_0007 <= (2**30)-1;
    i_distance_0008 <= (2**30)-1;
    i_distance_0009 <= (2**30)-1;
    i_distance_0010 <= (2**30)-1;
    i_distance_0011 <= (2**30)-1;
    i_distance_0012 <= (2**30)-1;
    i_distance_0013 <= (2**30)-1;
    i_distance_0014 <= (2**30)-1;
    i_distance_0015 <= (2**30)-1;
    i_distance_0016 <= (2**30)-1;
    i_distance_0017 <= (2**30)-1;
    i_distance_0018 <= (2**30)-1;
    i_distance_0019 <= (2**30)-1;
    i_distance_0020 <= (2**30)-1;
    i_distance_0021 <= (2**30)-1;
    i_distance_0022 <= (2**30)-1;
    i_distance_0023 <= (2**30)-1;
    i_distance_0024 <= (2**30)-1;
    i_distance_0025 <= (2**30)-1;
    i_distance_0026 <= (2**30)-1;
    i_distance_0027 <= (2**30)-1;
    i_distance_0028 <= (2**30)-1;
    i_distance_0029 <= (2**30)-1;
    i_distance_0030 <= (2**30)-1;
    i_distance_0031 <= (2**30)-1;
    i_distance_0032 <= (2**30)-1;
    i_distance_0033 <= (2**30)-1;
    i_distance_0034 <= (2**30)-1;
    i_distance_0035 <= (2**30)-1;
    i_distance_0036 <= (2**30)-1;
    i_distance_0037 <= (2**30)-1;
    i_distance_0038 <= (2**30)-1;
    i_distance_0039 <= (2**30)-1;
    i_distance_0040 <= (2**30)-1;
    i_distance_0041 <= (2**30)-1;
    i_distance_0042 <= (2**30)-1;
    i_distance_0043 <= (2**30)-1;
    i_distance_0044 <= (2**30)-1;
    i_distance_0045 <= (2**30)-1;
    i_distance_0046 <= (2**30)-1;
    i_distance_0047 <= (2**30)-1;
    i_distance_0048 <= (2**30)-1;
    i_distance_0049 <= (2**30)-1;
    i_distance_0050 <= (2**30)-1;
    i_distance_0051 <= (2**30)-1;
    i_distance_0052 <= (2**30)-1;
    i_distance_0053 <= (2**30)-1;
    i_distance_0054 <= (2**30)-1;
    i_distance_0055 <= (2**30)-1;
    i_distance_0056 <= (2**30)-1;
    i_distance_0057 <= (2**30)-1;
    i_distance_0058 <= (2**30)-1;
    i_distance_0059 <= (2**30)-1;
    i_distance_0060 <= (2**30)-1;
    i_distance_0061 <= (2**30)-1;
    i_distance_0062 <= (2**30)-1;
    i_distance_0063 <= (2**30)-1;
    correct_answer <= (2**30)-1;
    sync_wait_rising(clk, 10);
    rst <= not rst;
    sync_wait_rising(clk, 10);
    
    i_distance_0000 <= 588032;
    i_distance_0001 <= 4225;
    i_distance_0002 <= 12033;
    i_distance_0003 <= 3971;
    i_distance_0004 <= 212865;
    i_distance_0005 <= 996101;
    i_distance_0006 <= 1025922;
    i_distance_0007 <= 770950;
    i_distance_0008 <= 526214;
    i_distance_0009 <= 583689;
    i_distance_0010 <= 681609;
    i_distance_0011 <= 964621;
    i_distance_0012 <= 691605;
    i_distance_0013 <= 318486;
    i_distance_0014 <= 865303;
    i_distance_0015 <= 504855;
    i_distance_0016 <= 958358;
    i_distance_0017 <= 312858;
    i_distance_0018 <= 767259;
    i_distance_0019 <= 432539;
    i_distance_0020 <= 258462;
    i_distance_0021 <= 523556;
    i_distance_0022 <= 801191;
    i_distance_0023 <= 538538;
    i_distance_0024 <= 359341;
    i_distance_0025 <= 623022;
    i_distance_0026 <= 891445;
    i_distance_0027 <= 33846;
    i_distance_0028 <= 485817;
    i_distance_0029 <= 371131;
    i_distance_0030 <= 169276;
    i_distance_0031 <= 663230;
    i_distance_0032 <= 168895;
    i_distance_0033 <= 349377;
    i_distance_0034 <= 482881;
    i_distance_0035 <= 754625;
    i_distance_0036 <= 613699;
    i_distance_0037 <= 766792;
    i_distance_0038 <= 217675;
    i_distance_0039 <= 611020;
    i_distance_0040 <= 806732;
    i_distance_0041 <= 438221;
    i_distance_0042 <= 490316;
    i_distance_0043 <= 141134;
    i_distance_0044 <= 499282;
    i_distance_0045 <= 1023187;
    i_distance_0046 <= 887892;
    i_distance_0047 <= 160853;
    i_distance_0048 <= 887640;
    i_distance_0049 <= 964065;
    i_distance_0050 <= 338659;
    i_distance_0051 <= 15971;
    i_distance_0052 <= 495336;
    i_distance_0053 <= 865385;
    i_distance_0054 <= 588649;
    i_distance_0055 <= 601962;
    i_distance_0056 <= 691565;
    i_distance_0057 <= 403696;
    i_distance_0058 <= 973170;
    i_distance_0059 <= 243445;
    i_distance_0060 <= 206582;
    i_distance_0061 <= 327671;
    i_distance_0062 <= 241788;
    i_distance_0063 <= 814718;
    correct_answer <= 3971;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 622208;
    i_distance_0001 <= 51841;
    i_distance_0002 <= 614019;
    i_distance_0003 <= 185219;
    i_distance_0004 <= 482181;
    i_distance_0005 <= 271735;
    i_distance_0006 <= 1037701;
    i_distance_0007 <= 117768;
    i_distance_0008 <= 424972;
    i_distance_0009 <= 859149;
    i_distance_0010 <= 728977;
    i_distance_0011 <= 479890;
    i_distance_0012 <= 774549;
    i_distance_0013 <= 837144;
    i_distance_0014 <= 247576;
    i_distance_0015 <= 773659;
    i_distance_0016 <= 635163;
    i_distance_0017 <= 540321;
    i_distance_0018 <= 439678;
    i_distance_0019 <= 123171;
    i_distance_0020 <= 362281;
    i_distance_0021 <= 641710;
    i_distance_0022 <= 243249;
    i_distance_0023 <= 631731;
    i_distance_0024 <= 137013;
    i_distance_0025 <= 41781;
    i_distance_0026 <= 577848;
    i_distance_0027 <= 851768;
    i_distance_0028 <= 942781;
    i_distance_0029 <= 323008;
    i_distance_0030 <= 144193;
    i_distance_0031 <= 795200;
    i_distance_0032 <= 1028676;
    i_distance_0033 <= 356292;
    i_distance_0034 <= 986948;
    i_distance_0035 <= 185927;
    i_distance_0036 <= 433865;
    i_distance_0037 <= 110665;
    i_distance_0038 <= 564554;
    i_distance_0039 <= 874826;
    i_distance_0040 <= 897482;
    i_distance_0041 <= 10064;
    i_distance_0042 <= 170579;
    i_distance_0043 <= 584532;
    i_distance_0044 <= 702294;
    i_distance_0045 <= 99419;
    i_distance_0046 <= 368092;
    i_distance_0047 <= 556893;
    i_distance_0048 <= 211037;
    i_distance_0049 <= 801887;
    i_distance_0050 <= 959712;
    i_distance_0051 <= 926180;
    i_distance_0052 <= 635622;
    i_distance_0053 <= 516199;
    i_distance_0054 <= 235625;
    i_distance_0055 <= 420843;
    i_distance_0056 <= 173163;
    i_distance_0057 <= 885871;
    i_distance_0058 <= 891121;
    i_distance_0059 <= 447985;
    i_distance_0060 <= 371319;
    i_distance_0061 <= 277371;
    i_distance_0062 <= 759422;
    i_distance_0063 <= 1047423;
    correct_answer <= 10064;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 599042;
    i_distance_0001 <= 678020;
    i_distance_0002 <= 620422;
    i_distance_0003 <= 185478;
    i_distance_0004 <= 726920;
    i_distance_0005 <= 1002521;
    i_distance_0006 <= 697625;
    i_distance_0007 <= 1024283;
    i_distance_0008 <= 235163;
    i_distance_0009 <= 563738;
    i_distance_0010 <= 983585;
    i_distance_0011 <= 333182;
    i_distance_0012 <= 941864;
    i_distance_0013 <= 438830;
    i_distance_0014 <= 16430;
    i_distance_0015 <= 818480;
    i_distance_0016 <= 313137;
    i_distance_0017 <= 255409;
    i_distance_0018 <= 4528;
    i_distance_0019 <= 323636;
    i_distance_0020 <= 229941;
    i_distance_0021 <= 247860;
    i_distance_0022 <= 509625;
    i_distance_0023 <= 125497;
    i_distance_0024 <= 222652;
    i_distance_0025 <= 433341;
    i_distance_0026 <= 23228;
    i_distance_0027 <= 659391;
    i_distance_0028 <= 267969;
    i_distance_0029 <= 229192;
    i_distance_0030 <= 545480;
    i_distance_0031 <= 452425;
    i_distance_0032 <= 523467;
    i_distance_0033 <= 78157;
    i_distance_0034 <= 956878;
    i_distance_0035 <= 151885;
    i_distance_0036 <= 365136;
    i_distance_0037 <= 851668;
    i_distance_0038 <= 867928;
    i_distance_0039 <= 911576;
    i_distance_0040 <= 307547;
    i_distance_0041 <= 253405;
    i_distance_0042 <= 192094;
    i_distance_0043 <= 140511;
    i_distance_0044 <= 632543;
    i_distance_0045 <= 315618;
    i_distance_0046 <= 519778;
    i_distance_0047 <= 549988;
    i_distance_0048 <= 647650;
    i_distance_0049 <= 620004;
    i_distance_0050 <= 698087;
    i_distance_0051 <= 52962;
    i_distance_0052 <= 779114;
    i_distance_0053 <= 653803;
    i_distance_0054 <= 619755;
    i_distance_0055 <= 294762;
    i_distance_0056 <= 647666;
    i_distance_0057 <= 5236;
    i_distance_0058 <= 504950;
    i_distance_0059 <= 871671;
    i_distance_0060 <= 31737;
    i_distance_0061 <= 974845;
    i_distance_0062 <= 1039230;
    i_distance_0063 <= 80639;
    correct_answer <= 4528;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 418690;
    i_distance_0001 <= 584198;
    i_distance_0002 <= 944521;
    i_distance_0003 <= 228745;
    i_distance_0004 <= 226829;
    i_distance_0005 <= 354704;
    i_distance_0006 <= 144381;
    i_distance_0007 <= 299025;
    i_distance_0008 <= 8977;
    i_distance_0009 <= 328852;
    i_distance_0010 <= 1021205;
    i_distance_0011 <= 80536;
    i_distance_0012 <= 335001;
    i_distance_0013 <= 514072;
    i_distance_0014 <= 747293;
    i_distance_0015 <= 232734;
    i_distance_0016 <= 426399;
    i_distance_0017 <= 81440;
    i_distance_0018 <= 216735;
    i_distance_0019 <= 14967;
    i_distance_0020 <= 705194;
    i_distance_0021 <= 861739;
    i_distance_0022 <= 691376;
    i_distance_0023 <= 482423;
    i_distance_0024 <= 619065;
    i_distance_0025 <= 414780;
    i_distance_0026 <= 867900;
    i_distance_0027 <= 1029056;
    i_distance_0028 <= 162757;
    i_distance_0029 <= 724808;
    i_distance_0030 <= 253258;
    i_distance_0031 <= 532940;
    i_distance_0032 <= 575822;
    i_distance_0033 <= 28751;
    i_distance_0034 <= 384719;
    i_distance_0035 <= 598863;
    i_distance_0036 <= 436818;
    i_distance_0037 <= 770903;
    i_distance_0038 <= 220413;
    i_distance_0039 <= 986971;
    i_distance_0040 <= 475869;
    i_distance_0041 <= 173149;
    i_distance_0042 <= 179679;
    i_distance_0043 <= 184799;
    i_distance_0044 <= 507389;
    i_distance_0045 <= 744930;
    i_distance_0046 <= 641123;
    i_distance_0047 <= 576356;
    i_distance_0048 <= 839140;
    i_distance_0049 <= 462970;
    i_distance_0050 <= 631910;
    i_distance_0051 <= 1034466;
    i_distance_0052 <= 566891;
    i_distance_0053 <= 651118;
    i_distance_0054 <= 386289;
    i_distance_0055 <= 1014257;
    i_distance_0056 <= 84212;
    i_distance_0057 <= 406518;
    i_distance_0058 <= 544503;
    i_distance_0059 <= 932090;
    i_distance_0060 <= 439803;
    i_distance_0061 <= 845821;
    i_distance_0062 <= 990462;
    i_distance_0063 <= 946431;
    correct_answer <= 8977;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 125443;
    i_distance_0001 <= 690948;
    i_distance_0002 <= 519430;
    i_distance_0003 <= 64648;
    i_distance_0004 <= 917129;
    i_distance_0005 <= 469002;
    i_distance_0006 <= 505610;
    i_distance_0007 <= 21133;
    i_distance_0008 <= 709518;
    i_distance_0009 <= 984722;
    i_distance_0010 <= 1005200;
    i_distance_0011 <= 961809;
    i_distance_0012 <= 818065;
    i_distance_0013 <= 449427;
    i_distance_0014 <= 259348;
    i_distance_0015 <= 944532;
    i_distance_0016 <= 752918;
    i_distance_0017 <= 257686;
    i_distance_0018 <= 163736;
    i_distance_0019 <= 692632;
    i_distance_0020 <= 99605;
    i_distance_0021 <= 823320;
    i_distance_0022 <= 259228;
    i_distance_0023 <= 959645;
    i_distance_0024 <= 541;
    i_distance_0025 <= 820383;
    i_distance_0026 <= 1044895;
    i_distance_0027 <= 367643;
    i_distance_0028 <= 436386;
    i_distance_0029 <= 142749;
    i_distance_0030 <= 328484;
    i_distance_0031 <= 674471;
    i_distance_0032 <= 845865;
    i_distance_0033 <= 906153;
    i_distance_0034 <= 129453;
    i_distance_0035 <= 250547;
    i_distance_0036 <= 688699;
    i_distance_0037 <= 701883;
    i_distance_0038 <= 1026747;
    i_distance_0039 <= 579006;
    i_distance_0040 <= 508098;
    i_distance_0041 <= 274245;
    i_distance_0042 <= 560582;
    i_distance_0043 <= 107977;
    i_distance_0044 <= 40266;
    i_distance_0045 <= 428749;
    i_distance_0046 <= 1016400;
    i_distance_0047 <= 661715;
    i_distance_0048 <= 305366;
    i_distance_0049 <= 941278;
    i_distance_0050 <= 432993;
    i_distance_0051 <= 868066;
    i_distance_0052 <= 703841;
    i_distance_0053 <= 829669;
    i_distance_0054 <= 863742;
    i_distance_0055 <= 430950;
    i_distance_0056 <= 979434;
    i_distance_0057 <= 809964;
    i_distance_0058 <= 914287;
    i_distance_0059 <= 981873;
    i_distance_0060 <= 72441;
    i_distance_0061 <= 721658;
    i_distance_0062 <= 1026427;
    i_distance_0063 <= 315262;
    correct_answer <= 541;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 782208;
    i_distance_0001 <= 131843;
    i_distance_0002 <= 688003;
    i_distance_0003 <= 81797;
    i_distance_0004 <= 602629;
    i_distance_0005 <= 1040646;
    i_distance_0006 <= 990084;
    i_distance_0007 <= 258830;
    i_distance_0008 <= 853903;
    i_distance_0009 <= 253968;
    i_distance_0010 <= 112529;
    i_distance_0011 <= 402961;
    i_distance_0012 <= 410128;
    i_distance_0013 <= 850710;
    i_distance_0014 <= 903288;
    i_distance_0015 <= 127388;
    i_distance_0016 <= 1034270;
    i_distance_0017 <= 676639;
    i_distance_0018 <= 825890;
    i_distance_0019 <= 13474;
    i_distance_0020 <= 787491;
    i_distance_0021 <= 222249;
    i_distance_0022 <= 732206;
    i_distance_0023 <= 704303;
    i_distance_0024 <= 352817;
    i_distance_0025 <= 743604;
    i_distance_0026 <= 661687;
    i_distance_0027 <= 849722;
    i_distance_0028 <= 448320;
    i_distance_0029 <= 785090;
    i_distance_0030 <= 421315;
    i_distance_0031 <= 340674;
    i_distance_0032 <= 332485;
    i_distance_0033 <= 252742;
    i_distance_0034 <= 658503;
    i_distance_0035 <= 435016;
    i_distance_0036 <= 1018692;
    i_distance_0037 <= 161610;
    i_distance_0038 <= 778572;
    i_distance_0039 <= 175826;
    i_distance_0040 <= 765139;
    i_distance_0041 <= 118488;
    i_distance_0042 <= 139355;
    i_distance_0043 <= 1025116;
    i_distance_0044 <= 737884;
    i_distance_0045 <= 1048027;
    i_distance_0046 <= 876513;
    i_distance_0047 <= 836071;
    i_distance_0048 <= 575080;
    i_distance_0049 <= 732648;
    i_distance_0050 <= 861168;
    i_distance_0051 <= 875248;
    i_distance_0052 <= 682994;
    i_distance_0053 <= 790258;
    i_distance_0054 <= 418803;
    i_distance_0055 <= 538613;
    i_distance_0056 <= 791798;
    i_distance_0057 <= 812151;
    i_distance_0058 <= 323960;
    i_distance_0059 <= 710386;
    i_distance_0060 <= 752762;
    i_distance_0061 <= 377331;
    i_distance_0062 <= 530685;
    i_distance_0063 <= 671103;
    correct_answer <= 13474;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 795392;
    i_distance_0001 <= 44801;
    i_distance_0002 <= 156931;
    i_distance_0003 <= 284549;
    i_distance_0004 <= 880904;
    i_distance_0005 <= 805258;
    i_distance_0006 <= 857230;
    i_distance_0007 <= 638607;
    i_distance_0008 <= 382228;
    i_distance_0009 <= 848277;
    i_distance_0010 <= 319510;
    i_distance_0011 <= 350491;
    i_distance_0012 <= 523549;
    i_distance_0013 <= 918941;
    i_distance_0014 <= 557088;
    i_distance_0015 <= 963745;
    i_distance_0016 <= 372256;
    i_distance_0017 <= 281637;
    i_distance_0018 <= 373158;
    i_distance_0019 <= 167973;
    i_distance_0020 <= 172198;
    i_distance_0021 <= 816552;
    i_distance_0022 <= 608170;
    i_distance_0023 <= 324523;
    i_distance_0024 <= 143403;
    i_distance_0025 <= 667819;
    i_distance_0026 <= 512684;
    i_distance_0027 <= 313387;
    i_distance_0028 <= 1032624;
    i_distance_0029 <= 565937;
    i_distance_0030 <= 66865;
    i_distance_0031 <= 898604;
    i_distance_0032 <= 317101;
    i_distance_0033 <= 684479;
    i_distance_0034 <= 235585;
    i_distance_0035 <= 729794;
    i_distance_0036 <= 917441;
    i_distance_0037 <= 722756;
    i_distance_0038 <= 1022917;
    i_distance_0039 <= 256966;
    i_distance_0040 <= 748871;
    i_distance_0041 <= 600648;
    i_distance_0042 <= 735046;
    i_distance_0043 <= 407375;
    i_distance_0044 <= 567124;
    i_distance_0045 <= 918743;
    i_distance_0046 <= 460378;
    i_distance_0047 <= 244060;
    i_distance_0048 <= 579037;
    i_distance_0049 <= 318940;
    i_distance_0050 <= 795620;
    i_distance_0051 <= 548070;
    i_distance_0052 <= 226151;
    i_distance_0053 <= 903146;
    i_distance_0054 <= 214891;
    i_distance_0055 <= 161190;
    i_distance_0056 <= 954733;
    i_distance_0057 <= 707440;
    i_distance_0058 <= 529906;
    i_distance_0059 <= 665846;
    i_distance_0060 <= 503287;
    i_distance_0061 <= 1021944;
    i_distance_0062 <= 418940;
    i_distance_0063 <= 814205;
    correct_answer <= 44801;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 1022724;
    i_distance_0001 <= 520073;
    i_distance_0002 <= 996106;
    i_distance_0003 <= 273802;
    i_distance_0004 <= 727691;
    i_distance_0005 <= 493067;
    i_distance_0006 <= 605710;
    i_distance_0007 <= 806541;
    i_distance_0008 <= 548747;
    i_distance_0009 <= 81425;
    i_distance_0010 <= 395026;
    i_distance_0011 <= 830231;
    i_distance_0012 <= 1014808;
    i_distance_0013 <= 656281;
    i_distance_0014 <= 386202;
    i_distance_0015 <= 743581;
    i_distance_0016 <= 157854;
    i_distance_0017 <= 805534;
    i_distance_0018 <= 628518;
    i_distance_0019 <= 661671;
    i_distance_0020 <= 133031;
    i_distance_0021 <= 921000;
    i_distance_0022 <= 477613;
    i_distance_0023 <= 781231;
    i_distance_0024 <= 871733;
    i_distance_0025 <= 562489;
    i_distance_0026 <= 942652;
    i_distance_0027 <= 671167;
    i_distance_0028 <= 622022;
    i_distance_0029 <= 202697;
    i_distance_0030 <= 225225;
    i_distance_0031 <= 94154;
    i_distance_0032 <= 763724;
    i_distance_0033 <= 399309;
    i_distance_0034 <= 726222;
    i_distance_0035 <= 463183;
    i_distance_0036 <= 873167;
    i_distance_0037 <= 18383;
    i_distance_0038 <= 799568;
    i_distance_0039 <= 318291;
    i_distance_0040 <= 279896;
    i_distance_0041 <= 413656;
    i_distance_0042 <= 661339;
    i_distance_0043 <= 188507;
    i_distance_0044 <= 470875;
    i_distance_0045 <= 907998;
    i_distance_0046 <= 69343;
    i_distance_0047 <= 1025889;
    i_distance_0048 <= 79970;
    i_distance_0049 <= 491878;
    i_distance_0050 <= 656744;
    i_distance_0051 <= 151273;
    i_distance_0052 <= 761964;
    i_distance_0053 <= 63854;
    i_distance_0054 <= 866799;
    i_distance_0055 <= 761326;
    i_distance_0056 <= 828915;
    i_distance_0057 <= 750964;
    i_distance_0058 <= 1034485;
    i_distance_0059 <= 267764;
    i_distance_0060 <= 894711;
    i_distance_0061 <= 628469;
    i_distance_0062 <= 760950;
    i_distance_0063 <= 533886;
    correct_answer <= 18383;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 694787;
    i_distance_0001 <= 12934;
    i_distance_0002 <= 75399;
    i_distance_0003 <= 375432;
    i_distance_0004 <= 664073;
    i_distance_0005 <= 101774;
    i_distance_0006 <= 430863;
    i_distance_0007 <= 747408;
    i_distance_0008 <= 235026;
    i_distance_0009 <= 1011476;
    i_distance_0010 <= 541722;
    i_distance_0011 <= 480796;
    i_distance_0012 <= 963229;
    i_distance_0013 <= 13820;
    i_distance_0014 <= 26790;
    i_distance_0015 <= 287527;
    i_distance_0016 <= 84647;
    i_distance_0017 <= 564905;
    i_distance_0018 <= 193066;
    i_distance_0019 <= 580652;
    i_distance_0020 <= 292269;
    i_distance_0021 <= 144813;
    i_distance_0022 <= 971950;
    i_distance_0023 <= 139183;
    i_distance_0024 <= 621233;
    i_distance_0025 <= 872881;
    i_distance_0026 <= 497076;
    i_distance_0027 <= 226232;
    i_distance_0028 <= 850233;
    i_distance_0029 <= 177209;
    i_distance_0030 <= 161723;
    i_distance_0031 <= 190012;
    i_distance_0032 <= 675643;
    i_distance_0033 <= 119996;
    i_distance_0034 <= 818367;
    i_distance_0035 <= 838084;
    i_distance_0036 <= 909638;
    i_distance_0037 <= 543049;
    i_distance_0038 <= 38732;
    i_distance_0039 <= 708687;
    i_distance_0040 <= 607055;
    i_distance_0041 <= 348241;
    i_distance_0042 <= 995922;
    i_distance_0043 <= 267087;
    i_distance_0044 <= 467157;
    i_distance_0045 <= 467029;
    i_distance_0046 <= 798683;
    i_distance_0047 <= 27485;
    i_distance_0048 <= 277472;
    i_distance_0049 <= 130789;
    i_distance_0050 <= 1021925;
    i_distance_0051 <= 245095;
    i_distance_0052 <= 73469;
    i_distance_0053 <= 567402;
    i_distance_0054 <= 622313;
    i_distance_0055 <= 25208;
    i_distance_0056 <= 305132;
    i_distance_0057 <= 609134;
    i_distance_0058 <= 658928;
    i_distance_0059 <= 928882;
    i_distance_0060 <= 144248;
    i_distance_0061 <= 288378;
    i_distance_0062 <= 889212;
    i_distance_0063 <= 731901;
    correct_answer <= 12934;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 509186;
    i_distance_0001 <= 809220;
    i_distance_0002 <= 301700;
    i_distance_0003 <= 871816;
    i_distance_0004 <= 401547;
    i_distance_0005 <= 1041681;
    i_distance_0006 <= 1002393;
    i_distance_0007 <= 911258;
    i_distance_0008 <= 623388;
    i_distance_0009 <= 143005;
    i_distance_0010 <= 326814;
    i_distance_0011 <= 888607;
    i_distance_0012 <= 492959;
    i_distance_0013 <= 88476;
    i_distance_0014 <= 441886;
    i_distance_0015 <= 61853;
    i_distance_0016 <= 588833;
    i_distance_0017 <= 244899;
    i_distance_0018 <= 920742;
    i_distance_0019 <= 740902;
    i_distance_0020 <= 708011;
    i_distance_0021 <= 44459;
    i_distance_0022 <= 674605;
    i_distance_0023 <= 182318;
    i_distance_0024 <= 724017;
    i_distance_0025 <= 95282;
    i_distance_0026 <= 951860;
    i_distance_0027 <= 338613;
    i_distance_0028 <= 1047860;
    i_distance_0029 <= 156087;
    i_distance_0030 <= 548279;
    i_distance_0031 <= 190266;
    i_distance_0032 <= 634172;
    i_distance_0033 <= 948415;
    i_distance_0034 <= 860224;
    i_distance_0035 <= 174656;
    i_distance_0036 <= 825536;
    i_distance_0037 <= 19523;
    i_distance_0038 <= 671551;
    i_distance_0039 <= 466630;
    i_distance_0040 <= 207051;
    i_distance_0041 <= 378445;
    i_distance_0042 <= 956111;
    i_distance_0043 <= 929616;
    i_distance_0044 <= 148433;
    i_distance_0045 <= 968143;
    i_distance_0046 <= 913877;
    i_distance_0047 <= 263894;
    i_distance_0048 <= 413534;
    i_distance_0049 <= 634081;
    i_distance_0050 <= 799844;
    i_distance_0051 <= 746854;
    i_distance_0052 <= 583146;
    i_distance_0053 <= 676588;
    i_distance_0054 <= 3183;
    i_distance_0055 <= 574960;
    i_distance_0056 <= 303219;
    i_distance_0057 <= 712822;
    i_distance_0058 <= 263031;
    i_distance_0059 <= 1021433;
    i_distance_0060 <= 705274;
    i_distance_0061 <= 542972;
    i_distance_0062 <= 967165;
    i_distance_0063 <= 357630;
    correct_answer <= 3183;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 912769;
    i_distance_0001 <= 514306;
    i_distance_0002 <= 225924;
    i_distance_0003 <= 267141;
    i_distance_0004 <= 648838;
    i_distance_0005 <= 986887;
    i_distance_0006 <= 100488;
    i_distance_0007 <= 713991;
    i_distance_0008 <= 142869;
    i_distance_0009 <= 72855;
    i_distance_0010 <= 202521;
    i_distance_0011 <= 912026;
    i_distance_0012 <= 680347;
    i_distance_0013 <= 94620;
    i_distance_0014 <= 163609;
    i_distance_0015 <= 683806;
    i_distance_0016 <= 640671;
    i_distance_0017 <= 38432;
    i_distance_0018 <= 965282;
    i_distance_0019 <= 466342;
    i_distance_0020 <= 927912;
    i_distance_0021 <= 22570;
    i_distance_0022 <= 604588;
    i_distance_0023 <= 446384;
    i_distance_0024 <= 822576;
    i_distance_0025 <= 738356;
    i_distance_0026 <= 112311;
    i_distance_0027 <= 846651;
    i_distance_0028 <= 341819;
    i_distance_0029 <= 1001660;
    i_distance_0030 <= 3262;
    i_distance_0031 <= 148928;
    i_distance_0032 <= 995265;
    i_distance_0033 <= 472643;
    i_distance_0034 <= 544711;
    i_distance_0035 <= 964942;
    i_distance_0036 <= 480594;
    i_distance_0037 <= 290899;
    i_distance_0038 <= 204919;
    i_distance_0039 <= 583769;
    i_distance_0040 <= 304986;
    i_distance_0041 <= 816987;
    i_distance_0042 <= 546267;
    i_distance_0043 <= 478429;
    i_distance_0044 <= 41566;
    i_distance_0045 <= 23776;
    i_distance_0046 <= 1026528;
    i_distance_0047 <= 760162;
    i_distance_0048 <= 763491;
    i_distance_0049 <= 558818;
    i_distance_0050 <= 1019111;
    i_distance_0051 <= 188908;
    i_distance_0052 <= 972016;
    i_distance_0053 <= 235505;
    i_distance_0054 <= 302450;
    i_distance_0055 <= 670194;
    i_distance_0056 <= 449523;
    i_distance_0057 <= 967926;
    i_distance_0058 <= 18935;
    i_distance_0059 <= 24952;
    i_distance_0060 <= 207222;
    i_distance_0061 <= 369659;
    i_distance_0062 <= 153853;
    i_distance_0063 <= 476671;
    correct_answer <= 3262;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 780928;
    i_distance_0001 <= 378370;
    i_distance_0002 <= 452738;
    i_distance_0003 <= 825091;
    i_distance_0004 <= 277255;
    i_distance_0005 <= 958216;
    i_distance_0006 <= 254217;
    i_distance_0007 <= 326666;
    i_distance_0008 <= 868106;
    i_distance_0009 <= 605835;
    i_distance_0010 <= 675976;
    i_distance_0011 <= 273930;
    i_distance_0012 <= 860297;
    i_distance_0013 <= 183568;
    i_distance_0014 <= 821267;
    i_distance_0015 <= 141593;
    i_distance_0016 <= 757914;
    i_distance_0017 <= 241947;
    i_distance_0018 <= 1019804;
    i_distance_0019 <= 771354;
    i_distance_0020 <= 970399;
    i_distance_0021 <= 571296;
    i_distance_0022 <= 889631;
    i_distance_0023 <= 1442;
    i_distance_0024 <= 181922;
    i_distance_0025 <= 121122;
    i_distance_0026 <= 368429;
    i_distance_0027 <= 352048;
    i_distance_0028 <= 187313;
    i_distance_0029 <= 518833;
    i_distance_0030 <= 541360;
    i_distance_0031 <= 630580;
    i_distance_0032 <= 276662;
    i_distance_0033 <= 549816;
    i_distance_0034 <= 856889;
    i_distance_0035 <= 299454;
    i_distance_0036 <= 180799;
    i_distance_0037 <= 856129;
    i_distance_0038 <= 797635;
    i_distance_0039 <= 10820;
    i_distance_0040 <= 272072;
    i_distance_0041 <= 283724;
    i_distance_0042 <= 215760;
    i_distance_0043 <= 425938;
    i_distance_0044 <= 239828;
    i_distance_0045 <= 444245;
    i_distance_0046 <= 843481;
    i_distance_0047 <= 1018841;
    i_distance_0048 <= 293980;
    i_distance_0049 <= 946653;
    i_distance_0050 <= 665825;
    i_distance_0051 <= 758754;
    i_distance_0052 <= 406882;
    i_distance_0053 <= 210661;
    i_distance_0054 <= 412134;
    i_distance_0055 <= 66152;
    i_distance_0056 <= 269545;
    i_distance_0057 <= 92008;
    i_distance_0058 <= 646510;
    i_distance_0059 <= 151026;
    i_distance_0060 <= 490740;
    i_distance_0061 <= 419063;
    i_distance_0062 <= 454265;
    i_distance_0063 <= 748287;
    correct_answer <= 1442;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 627072;
    i_distance_0001 <= 913025;
    i_distance_0002 <= 885892;
    i_distance_0003 <= 664457;
    i_distance_0004 <= 359948;
    i_distance_0005 <= 806029;
    i_distance_0006 <= 505358;
    i_distance_0007 <= 709268;
    i_distance_0008 <= 130070;
    i_distance_0009 <= 14103;
    i_distance_0010 <= 418842;
    i_distance_0011 <= 2716;
    i_distance_0012 <= 44828;
    i_distance_0013 <= 38047;
    i_distance_0014 <= 651424;
    i_distance_0015 <= 980258;
    i_distance_0016 <= 921635;
    i_distance_0017 <= 290341;
    i_distance_0018 <= 327721;
    i_distance_0019 <= 610094;
    i_distance_0020 <= 284081;
    i_distance_0021 <= 79160;
    i_distance_0022 <= 753080;
    i_distance_0023 <= 391294;
    i_distance_0024 <= 636224;
    i_distance_0025 <= 693443;
    i_distance_0026 <= 24644;
    i_distance_0027 <= 1027783;
    i_distance_0028 <= 666440;
    i_distance_0029 <= 844362;
    i_distance_0030 <= 941771;
    i_distance_0031 <= 415051;
    i_distance_0032 <= 659021;
    i_distance_0033 <= 900042;
    i_distance_0034 <= 46803;
    i_distance_0035 <= 938964;
    i_distance_0036 <= 428501;
    i_distance_0037 <= 249557;
    i_distance_0038 <= 45397;
    i_distance_0039 <= 616792;
    i_distance_0040 <= 446425;
    i_distance_0041 <= 949374;
    i_distance_0042 <= 334298;
    i_distance_0043 <= 380635;
    i_distance_0044 <= 157151;
    i_distance_0045 <= 896992;
    i_distance_0046 <= 608994;
    i_distance_0047 <= 132835;
    i_distance_0048 <= 372068;
    i_distance_0049 <= 645734;
    i_distance_0050 <= 666982;
    i_distance_0051 <= 714347;
    i_distance_0052 <= 854123;
    i_distance_0053 <= 310125;
    i_distance_0054 <= 957807;
    i_distance_0055 <= 922865;
    i_distance_0056 <= 624883;
    i_distance_0057 <= 861811;
    i_distance_0058 <= 231029;
    i_distance_0059 <= 271734;
    i_distance_0060 <= 614903;
    i_distance_0061 <= 258934;
    i_distance_0062 <= 716669;
    i_distance_0063 <= 1046782;
    correct_answer <= 2716;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 779385;
    i_distance_0001 <= 669188;
    i_distance_0002 <= 735108;
    i_distance_0003 <= 650122;
    i_distance_0004 <= 370296;
    i_distance_0005 <= 569100;
    i_distance_0006 <= 584718;
    i_distance_0007 <= 972943;
    i_distance_0008 <= 29839;
    i_distance_0009 <= 491026;
    i_distance_0010 <= 160403;
    i_distance_0011 <= 85525;
    i_distance_0012 <= 772248;
    i_distance_0013 <= 1028252;
    i_distance_0014 <= 727709;
    i_distance_0015 <= 828191;
    i_distance_0016 <= 823845;
    i_distance_0017 <= 383141;
    i_distance_0018 <= 293032;
    i_distance_0019 <= 773802;
    i_distance_0020 <= 36395;
    i_distance_0021 <= 712874;
    i_distance_0022 <= 345902;
    i_distance_0023 <= 539695;
    i_distance_0024 <= 198319;
    i_distance_0025 <= 397617;
    i_distance_0026 <= 530484;
    i_distance_0027 <= 604725;
    i_distance_0028 <= 102198;
    i_distance_0029 <= 34871;
    i_distance_0030 <= 277176;
    i_distance_0031 <= 369337;
    i_distance_0032 <= 37689;
    i_distance_0033 <= 589116;
    i_distance_0034 <= 278079;
    i_distance_0035 <= 100288;
    i_distance_0036 <= 340417;
    i_distance_0037 <= 317503;
    i_distance_0038 <= 231492;
    i_distance_0039 <= 459335;
    i_distance_0040 <= 838344;
    i_distance_0041 <= 762444;
    i_distance_0042 <= 133582;
    i_distance_0043 <= 836303;
    i_distance_0044 <= 221264;
    i_distance_0045 <= 265426;
    i_distance_0046 <= 656596;
    i_distance_0047 <= 1023832;
    i_distance_0048 <= 752985;
    i_distance_0049 <= 695130;
    i_distance_0050 <= 839645;
    i_distance_0051 <= 320863;
    i_distance_0052 <= 781664;
    i_distance_0053 <= 234847;
    i_distance_0054 <= 465384;
    i_distance_0055 <= 229993;
    i_distance_0056 <= 412141;
    i_distance_0057 <= 983277;
    i_distance_0058 <= 994804;
    i_distance_0059 <= 304502;
    i_distance_0060 <= 867447;
    i_distance_0061 <= 819576;
    i_distance_0062 <= 827766;
    i_distance_0063 <= 535549;
    correct_answer <= 29839;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 445184;
    i_distance_0001 <= 736768;
    i_distance_0002 <= 889730;
    i_distance_0003 <= 1004420;
    i_distance_0004 <= 400132;
    i_distance_0005 <= 122888;
    i_distance_0006 <= 65674;
    i_distance_0007 <= 512140;
    i_distance_0008 <= 159247;
    i_distance_0009 <= 396049;
    i_distance_0010 <= 816145;
    i_distance_0011 <= 136979;
    i_distance_0012 <= 72980;
    i_distance_0013 <= 7840;
    i_distance_0014 <= 756897;
    i_distance_0015 <= 779299;
    i_distance_0016 <= 859556;
    i_distance_0017 <= 197412;
    i_distance_0018 <= 459044;
    i_distance_0019 <= 287145;
    i_distance_0020 <= 803754;
    i_distance_0021 <= 502698;
    i_distance_0022 <= 514474;
    i_distance_0023 <= 974765;
    i_distance_0024 <= 879659;
    i_distance_0025 <= 722990;
    i_distance_0026 <= 583605;
    i_distance_0027 <= 361142;
    i_distance_0028 <= 769591;
    i_distance_0029 <= 470327;
    i_distance_0030 <= 138299;
    i_distance_0031 <= 452671;
    i_distance_0032 <= 729409;
    i_distance_0033 <= 794308;
    i_distance_0034 <= 347718;
    i_distance_0035 <= 33095;
    i_distance_0036 <= 51528;
    i_distance_0037 <= 889415;
    i_distance_0038 <= 44493;
    i_distance_0039 <= 493647;
    i_distance_0040 <= 48213;
    i_distance_0041 <= 500694;
    i_distance_0042 <= 585173;
    i_distance_0043 <= 272984;
    i_distance_0044 <= 360793;
    i_distance_0045 <= 830677;
    i_distance_0046 <= 160219;
    i_distance_0047 <= 952667;
    i_distance_0048 <= 319454;
    i_distance_0049 <= 176351;
    i_distance_0050 <= 413797;
    i_distance_0051 <= 762213;
    i_distance_0052 <= 554985;
    i_distance_0053 <= 573035;
    i_distance_0054 <= 253547;
    i_distance_0055 <= 46189;
    i_distance_0056 <= 695149;
    i_distance_0057 <= 284527;
    i_distance_0058 <= 969199;
    i_distance_0059 <= 89461;
    i_distance_0060 <= 466934;
    i_distance_0061 <= 863738;
    i_distance_0062 <= 449790;
    i_distance_0063 <= 152447;
    correct_answer <= 7840;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 170497;
    i_distance_0001 <= 466306;
    i_distance_0002 <= 668678;
    i_distance_0003 <= 669453;
    i_distance_0004 <= 814477;
    i_distance_0005 <= 1024525;
    i_distance_0006 <= 434957;
    i_distance_0007 <= 415382;
    i_distance_0008 <= 957846;
    i_distance_0009 <= 689942;
    i_distance_0010 <= 214678;
    i_distance_0011 <= 971419;
    i_distance_0012 <= 115868;
    i_distance_0013 <= 422942;
    i_distance_0014 <= 912288;
    i_distance_0015 <= 713123;
    i_distance_0016 <= 289955;
    i_distance_0017 <= 534951;
    i_distance_0018 <= 317735;
    i_distance_0019 <= 437931;
    i_distance_0020 <= 328749;
    i_distance_0021 <= 798260;
    i_distance_0022 <= 438072;
    i_distance_0023 <= 398904;
    i_distance_0024 <= 1030458;
    i_distance_0025 <= 97853;
    i_distance_0026 <= 885310;
    i_distance_0027 <= 543807;
    i_distance_0028 <= 1040576;
    i_distance_0029 <= 103289;
    i_distance_0030 <= 48969;
    i_distance_0031 <= 279370;
    i_distance_0032 <= 539466;
    i_distance_0033 <= 117066;
    i_distance_0034 <= 255436;
    i_distance_0035 <= 747982;
    i_distance_0036 <= 227786;
    i_distance_0037 <= 1028553;
    i_distance_0038 <= 978513;
    i_distance_0039 <= 204618;
    i_distance_0040 <= 751315;
    i_distance_0041 <= 324692;
    i_distance_0042 <= 725461;
    i_distance_0043 <= 266838;
    i_distance_0044 <= 37333;
    i_distance_0045 <= 46296;
    i_distance_0046 <= 461918;
    i_distance_0047 <= 775392;
    i_distance_0048 <= 901474;
    i_distance_0049 <= 45026;
    i_distance_0050 <= 766820;
    i_distance_0051 <= 964324;
    i_distance_0052 <= 411235;
    i_distance_0053 <= 591079;
    i_distance_0054 <= 654563;
    i_distance_0055 <= 572009;
    i_distance_0056 <= 980714;
    i_distance_0057 <= 466924;
    i_distance_0058 <= 312686;
    i_distance_0059 <= 816495;
    i_distance_0060 <= 1033331;
    i_distance_0061 <= 886774;
    i_distance_0062 <= 548089;
    i_distance_0063 <= 78716;
    correct_answer <= 37333;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 385540;
    i_distance_0001 <= 130310;
    i_distance_0002 <= 251655;
    i_distance_0003 <= 730631;
    i_distance_0004 <= 382729;
    i_distance_0005 <= 269577;
    i_distance_0006 <= 452875;
    i_distance_0007 <= 803340;
    i_distance_0008 <= 623117;
    i_distance_0009 <= 847502;
    i_distance_0010 <= 974478;
    i_distance_0011 <= 436238;
    i_distance_0012 <= 166033;
    i_distance_0013 <= 274581;
    i_distance_0014 <= 315163;
    i_distance_0015 <= 274077;
    i_distance_0016 <= 181151;
    i_distance_0017 <= 447393;
    i_distance_0018 <= 559393;
    i_distance_0019 <= 797858;
    i_distance_0020 <= 125862;
    i_distance_0021 <= 24488;
    i_distance_0022 <= 657578;
    i_distance_0023 <= 948651;
    i_distance_0024 <= 173869;
    i_distance_0025 <= 601006;
    i_distance_0026 <= 913969;
    i_distance_0027 <= 609202;
    i_distance_0028 <= 254514;
    i_distance_0029 <= 969652;
    i_distance_0030 <= 37682;
    i_distance_0031 <= 801078;
    i_distance_0032 <= 38713;
    i_distance_0033 <= 902463;
    i_distance_0034 <= 693571;
    i_distance_0035 <= 948936;
    i_distance_0036 <= 500809;
    i_distance_0037 <= 454731;
    i_distance_0038 <= 525643;
    i_distance_0039 <= 779853;
    i_distance_0040 <= 126287;
    i_distance_0041 <= 700752;
    i_distance_0042 <= 717781;
    i_distance_0043 <= 298072;
    i_distance_0044 <= 827226;
    i_distance_0045 <= 86621;
    i_distance_0046 <= 98655;
    i_distance_0047 <= 527200;
    i_distance_0048 <= 303456;
    i_distance_0049 <= 873186;
    i_distance_0050 <= 115301;
    i_distance_0051 <= 237414;
    i_distance_0052 <= 573054;
    i_distance_0053 <= 680175;
    i_distance_0054 <= 618224;
    i_distance_0055 <= 743409;
    i_distance_0056 <= 524660;
    i_distance_0057 <= 959349;
    i_distance_0058 <= 773750;
    i_distance_0059 <= 876411;
    i_distance_0060 <= 249596;
    i_distance_0061 <= 476669;
    i_distance_0062 <= 895998;
    i_distance_0063 <= 370943;
    correct_answer <= 24488;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 680065;
    i_distance_0001 <= 588161;
    i_distance_0002 <= 427908;
    i_distance_0003 <= 545925;
    i_distance_0004 <= 888967;
    i_distance_0005 <= 858505;
    i_distance_0006 <= 258314;
    i_distance_0007 <= 641043;
    i_distance_0008 <= 429588;
    i_distance_0009 <= 538133;
    i_distance_0010 <= 983190;
    i_distance_0011 <= 266648;
    i_distance_0012 <= 525978;
    i_distance_0013 <= 886305;
    i_distance_0014 <= 700321;
    i_distance_0015 <= 374947;
    i_distance_0016 <= 546468;
    i_distance_0017 <= 658211;
    i_distance_0018 <= 281506;
    i_distance_0019 <= 7844;
    i_distance_0020 <= 163115;
    i_distance_0021 <= 208172;
    i_distance_0022 <= 66093;
    i_distance_0023 <= 1004972;
    i_distance_0024 <= 170927;
    i_distance_0025 <= 844464;
    i_distance_0026 <= 739889;
    i_distance_0027 <= 613297;
    i_distance_0028 <= 171059;
    i_distance_0029 <= 631342;
    i_distance_0030 <= 838325;
    i_distance_0031 <= 319798;
    i_distance_0032 <= 267575;
    i_distance_0033 <= 702391;
    i_distance_0034 <= 1031737;
    i_distance_0035 <= 751036;
    i_distance_0036 <= 308546;
    i_distance_0037 <= 404422;
    i_distance_0038 <= 822471;
    i_distance_0039 <= 559815;
    i_distance_0040 <= 551369;
    i_distance_0041 <= 977486;
    i_distance_0042 <= 480719;
    i_distance_0043 <= 525520;
    i_distance_0044 <= 142287;
    i_distance_0045 <= 1015253;
    i_distance_0046 <= 775893;
    i_distance_0047 <= 743385;
    i_distance_0048 <= 369627;
    i_distance_0049 <= 612446;
    i_distance_0050 <= 448352;
    i_distance_0051 <= 879458;
    i_distance_0052 <= 193379;
    i_distance_0053 <= 333796;
    i_distance_0054 <= 532072;
    i_distance_0055 <= 79208;
    i_distance_0056 <= 569322;
    i_distance_0057 <= 622059;
    i_distance_0058 <= 146412;
    i_distance_0059 <= 616044;
    i_distance_0060 <= 380403;
    i_distance_0061 <= 969460;
    i_distance_0062 <= 420597;
    i_distance_0063 <= 392570;
    correct_answer <= 7844;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 456833;
    i_distance_0001 <= 613890;
    i_distance_0002 <= 925955;
    i_distance_0003 <= 27139;
    i_distance_0004 <= 1047943;
    i_distance_0005 <= 832267;
    i_distance_0006 <= 18443;
    i_distance_0007 <= 575883;
    i_distance_0008 <= 318862;
    i_distance_0009 <= 319123;
    i_distance_0010 <= 562708;
    i_distance_0011 <= 321173;
    i_distance_0012 <= 659989;
    i_distance_0013 <= 881304;
    i_distance_0014 <= 183965;
    i_distance_0015 <= 490271;
    i_distance_0016 <= 216354;
    i_distance_0017 <= 495782;
    i_distance_0018 <= 915366;
    i_distance_0019 <= 679336;
    i_distance_0020 <= 340905;
    i_distance_0021 <= 695335;
    i_distance_0022 <= 580272;
    i_distance_0023 <= 590257;
    i_distance_0024 <= 222514;
    i_distance_0025 <= 237107;
    i_distance_0026 <= 921266;
    i_distance_0027 <= 866483;
    i_distance_0028 <= 501558;
    i_distance_0029 <= 596538;
    i_distance_0030 <= 172860;
    i_distance_0031 <= 487228;
    i_distance_0032 <= 904770;
    i_distance_0033 <= 600003;
    i_distance_0034 <= 829379;
    i_distance_0035 <= 922564;
    i_distance_0036 <= 1037126;
    i_distance_0037 <= 816200;
    i_distance_0038 <= 813642;
    i_distance_0039 <= 567627;
    i_distance_0040 <= 902730;
    i_distance_0041 <= 739408;
    i_distance_0042 <= 499411;
    i_distance_0043 <= 779605;
    i_distance_0044 <= 691286;
    i_distance_0045 <= 512600;
    i_distance_0046 <= 975065;
    i_distance_0047 <= 458969;
    i_distance_0048 <= 312154;
    i_distance_0049 <= 1010780;
    i_distance_0050 <= 485472;
    i_distance_0051 <= 351329;
    i_distance_0052 <= 697442;
    i_distance_0053 <= 636902;
    i_distance_0054 <= 690663;
    i_distance_0055 <= 465643;
    i_distance_0056 <= 616683;
    i_distance_0057 <= 123374;
    i_distance_0058 <= 510064;
    i_distance_0059 <= 1020273;
    i_distance_0060 <= 32629;
    i_distance_0061 <= 193911;
    i_distance_0062 <= 843387;
    i_distance_0063 <= 766204;
    correct_answer <= 18443;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 188547;
    i_distance_0001 <= 382983;
    i_distance_0002 <= 472586;
    i_distance_0003 <= 13963;
    i_distance_0004 <= 175500;
    i_distance_0005 <= 967183;
    i_distance_0006 <= 875413;
    i_distance_0007 <= 378136;
    i_distance_0008 <= 549912;
    i_distance_0009 <= 1033496;
    i_distance_0010 <= 31514;
    i_distance_0011 <= 146715;
    i_distance_0012 <= 214819;
    i_distance_0013 <= 741797;
    i_distance_0014 <= 148391;
    i_distance_0015 <= 702759;
    i_distance_0016 <= 686507;
    i_distance_0017 <= 354863;
    i_distance_0018 <= 25008;
    i_distance_0019 <= 444465;
    i_distance_0020 <= 889138;
    i_distance_0021 <= 46518;
    i_distance_0022 <= 250679;
    i_distance_0023 <= 576312;
    i_distance_0024 <= 220090;
    i_distance_0025 <= 973758;
    i_distance_0026 <= 110274;
    i_distance_0027 <= 514245;
    i_distance_0028 <= 503238;
    i_distance_0029 <= 771015;
    i_distance_0030 <= 163655;
    i_distance_0031 <= 809033;
    i_distance_0032 <= 697034;
    i_distance_0033 <= 463052;
    i_distance_0034 <= 500815;
    i_distance_0035 <= 302416;
    i_distance_0036 <= 160721;
    i_distance_0037 <= 623570;
    i_distance_0038 <= 15183;
    i_distance_0039 <= 401620;
    i_distance_0040 <= 515283;
    i_distance_0041 <= 342480;
    i_distance_0042 <= 912983;
    i_distance_0043 <= 505945;
    i_distance_0044 <= 724442;
    i_distance_0045 <= 105179;
    i_distance_0046 <= 781787;
    i_distance_0047 <= 259808;
    i_distance_0048 <= 113762;
    i_distance_0049 <= 638563;
    i_distance_0050 <= 1011944;
    i_distance_0051 <= 670573;
    i_distance_0052 <= 884974;
    i_distance_0053 <= 357997;
    i_distance_0054 <= 578416;
    i_distance_0055 <= 692462;
    i_distance_0056 <= 604018;
    i_distance_0057 <= 998132;
    i_distance_0058 <= 484340;
    i_distance_0059 <= 318838;
    i_distance_0060 <= 5241;
    i_distance_0061 <= 374266;
    i_distance_0062 <= 78459;
    i_distance_0063 <= 903295;
    correct_answer <= 5241;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 720128;
    i_distance_0001 <= 646275;
    i_distance_0002 <= 1040516;
    i_distance_0003 <= 582149;
    i_distance_0004 <= 237446;
    i_distance_0005 <= 110727;
    i_distance_0006 <= 12935;
    i_distance_0007 <= 860168;
    i_distance_0008 <= 341131;
    i_distance_0009 <= 686478;
    i_distance_0010 <= 839314;
    i_distance_0011 <= 534041;
    i_distance_0012 <= 929562;
    i_distance_0013 <= 574745;
    i_distance_0014 <= 316574;
    i_distance_0015 <= 485023;
    i_distance_0016 <= 459168;
    i_distance_0017 <= 723488;
    i_distance_0018 <= 629155;
    i_distance_0019 <= 78499;
    i_distance_0020 <= 1020195;
    i_distance_0021 <= 440742;
    i_distance_0022 <= 920487;
    i_distance_0023 <= 288677;
    i_distance_0024 <= 1013673;
    i_distance_0025 <= 919467;
    i_distance_0026 <= 810412;
    i_distance_0027 <= 1010221;
    i_distance_0028 <= 564396;
    i_distance_0029 <= 520753;
    i_distance_0030 <= 717235;
    i_distance_0031 <= 871862;
    i_distance_0032 <= 363959;
    i_distance_0033 <= 374071;
    i_distance_0034 <= 302393;
    i_distance_0035 <= 958393;
    i_distance_0036 <= 219192;
    i_distance_0037 <= 777406;
    i_distance_0038 <= 467905;
    i_distance_0039 <= 85187;
    i_distance_0040 <= 659396;
    i_distance_0041 <= 514372;
    i_distance_0042 <= 873415;
    i_distance_0043 <= 106311;
    i_distance_0044 <= 505672;
    i_distance_0045 <= 127061;
    i_distance_0046 <= 511447;
    i_distance_0047 <= 360536;
    i_distance_0048 <= 508119;
    i_distance_0049 <= 675418;
    i_distance_0050 <= 314849;
    i_distance_0051 <= 639713;
    i_distance_0052 <= 706787;
    i_distance_0053 <= 476774;
    i_distance_0054 <= 378857;
    i_distance_0055 <= 839916;
    i_distance_0056 <= 442988;
    i_distance_0057 <= 663532;
    i_distance_0058 <= 67055;
    i_distance_0059 <= 563692;
    i_distance_0060 <= 856943;
    i_distance_0061 <= 591219;
    i_distance_0062 <= 334198;
    i_distance_0063 <= 71807;
    correct_answer <= 12935;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 831878;
    i_distance_0001 <= 287366;
    i_distance_0002 <= 631549;
    i_distance_0003 <= 698251;
    i_distance_0004 <= 248716;
    i_distance_0005 <= 563086;
    i_distance_0006 <= 293519;
    i_distance_0007 <= 495252;
    i_distance_0008 <= 980629;
    i_distance_0009 <= 327701;
    i_distance_0010 <= 1012887;
    i_distance_0011 <= 51097;
    i_distance_0012 <= 1025689;
    i_distance_0013 <= 448539;
    i_distance_0014 <= 233244;
    i_distance_0015 <= 169889;
    i_distance_0016 <= 954401;
    i_distance_0017 <= 760355;
    i_distance_0018 <= 156449;
    i_distance_0019 <= 21285;
    i_distance_0020 <= 814509;
    i_distance_0021 <= 570159;
    i_distance_0022 <= 858160;
    i_distance_0023 <= 549297;
    i_distance_0024 <= 321330;
    i_distance_0025 <= 124850;
    i_distance_0026 <= 1004472;
    i_distance_0027 <= 183865;
    i_distance_0028 <= 828600;
    i_distance_0029 <= 499772;
    i_distance_0030 <= 1037630;
    i_distance_0031 <= 399298;
    i_distance_0032 <= 578758;
    i_distance_0033 <= 56648;
    i_distance_0034 <= 1010892;
    i_distance_0035 <= 468429;
    i_distance_0036 <= 835791;
    i_distance_0037 <= 329423;
    i_distance_0038 <= 376657;
    i_distance_0039 <= 905938;
    i_distance_0040 <= 808274;
    i_distance_0041 <= 14801;
    i_distance_0042 <= 619989;
    i_distance_0043 <= 664534;
    i_distance_0044 <= 665434;
    i_distance_0045 <= 689755;
    i_distance_0046 <= 943709;
    i_distance_0047 <= 936672;
    i_distance_0048 <= 564194;
    i_distance_0049 <= 534246;
    i_distance_0050 <= 297318;
    i_distance_0051 <= 145129;
    i_distance_0052 <= 496490;
    i_distance_0053 <= 830062;
    i_distance_0054 <= 376304;
    i_distance_0055 <= 866033;
    i_distance_0056 <= 925938;
    i_distance_0057 <= 876287;
    i_distance_0058 <= 49009;
    i_distance_0059 <= 265209;
    i_distance_0060 <= 663674;
    i_distance_0061 <= 596733;
    i_distance_0062 <= 503806;
    i_distance_0063 <= 401279;
    correct_answer <= 14801;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 983040;
    i_distance_0001 <= 267905;
    i_distance_0002 <= 934916;
    i_distance_0003 <= 1005452;
    i_distance_0004 <= 82069;
    i_distance_0005 <= 456597;
    i_distance_0006 <= 390685;
    i_distance_0007 <= 222368;
    i_distance_0008 <= 128161;
    i_distance_0009 <= 832290;
    i_distance_0010 <= 144933;
    i_distance_0011 <= 243109;
    i_distance_0012 <= 1040805;
    i_distance_0013 <= 483240;
    i_distance_0014 <= 327081;
    i_distance_0015 <= 684200;
    i_distance_0016 <= 997675;
    i_distance_0017 <= 510509;
    i_distance_0018 <= 799277;
    i_distance_0019 <= 559536;
    i_distance_0020 <= 450996;
    i_distance_0021 <= 414776;
    i_distance_0022 <= 624057;
    i_distance_0023 <= 826685;
    i_distance_0024 <= 72381;
    i_distance_0025 <= 355519;
    i_distance_0026 <= 411072;
    i_distance_0027 <= 104513;
    i_distance_0028 <= 954946;
    i_distance_0029 <= 75331;
    i_distance_0030 <= 430276;
    i_distance_0031 <= 421060;
    i_distance_0032 <= 87114;
    i_distance_0033 <= 485838;
    i_distance_0034 <= 542159;
    i_distance_0035 <= 40144;
    i_distance_0036 <= 961489;
    i_distance_0037 <= 405456;
    i_distance_0038 <= 452054;
    i_distance_0039 <= 470615;
    i_distance_0040 <= 380888;
    i_distance_0041 <= 815190;
    i_distance_0042 <= 787677;
    i_distance_0043 <= 250590;
    i_distance_0044 <= 105309;
    i_distance_0045 <= 447072;
    i_distance_0046 <= 60384;
    i_distance_0047 <= 1008228;
    i_distance_0048 <= 995813;
    i_distance_0049 <= 242021;
    i_distance_0050 <= 379622;
    i_distance_0051 <= 108137;
    i_distance_0052 <= 960490;
    i_distance_0053 <= 681709;
    i_distance_0054 <= 985841;
    i_distance_0055 <= 260978;
    i_distance_0056 <= 832755;
    i_distance_0057 <= 330227;
    i_distance_0058 <= 991346;
    i_distance_0059 <= 282359;
    i_distance_0060 <= 978299;
    i_distance_0061 <= 756861;
    i_distance_0062 <= 535678;
    i_distance_0063 <= 268799;
    correct_answer <= 40144;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 725634;
    i_distance_0001 <= 73218;
    i_distance_0002 <= 778631;
    i_distance_0003 <= 952074;
    i_distance_0004 <= 469514;
    i_distance_0005 <= 963598;
    i_distance_0006 <= 697359;
    i_distance_0007 <= 387728;
    i_distance_0008 <= 459663;
    i_distance_0009 <= 9230;
    i_distance_0010 <= 103316;
    i_distance_0011 <= 200085;
    i_distance_0012 <= 987286;
    i_distance_0013 <= 100244;
    i_distance_0014 <= 157716;
    i_distance_0015 <= 186776;
    i_distance_0016 <= 193178;
    i_distance_0017 <= 54171;
    i_distance_0018 <= 955930;
    i_distance_0019 <= 795037;
    i_distance_0020 <= 57635;
    i_distance_0021 <= 999846;
    i_distance_0022 <= 819622;
    i_distance_0023 <= 877864;
    i_distance_0024 <= 179497;
    i_distance_0025 <= 468266;
    i_distance_0026 <= 450988;
    i_distance_0027 <= 516269;
    i_distance_0028 <= 288429;
    i_distance_0029 <= 658351;
    i_distance_0030 <= 31532;
    i_distance_0031 <= 341169;
    i_distance_0032 <= 507058;
    i_distance_0033 <= 555053;
    i_distance_0034 <= 836020;
    i_distance_0035 <= 360119;
    i_distance_0036 <= 666553;
    i_distance_0037 <= 600637;
    i_distance_0038 <= 846013;
    i_distance_0039 <= 1009981;
    i_distance_0040 <= 284354;
    i_distance_0041 <= 322498;
    i_distance_0042 <= 723140;
    i_distance_0043 <= 244418;
    i_distance_0044 <= 131269;
    i_distance_0045 <= 1044040;
    i_distance_0046 <= 316235;
    i_distance_0047 <= 464849;
    i_distance_0048 <= 676434;
    i_distance_0049 <= 564055;
    i_distance_0050 <= 719195;
    i_distance_0051 <= 405852;
    i_distance_0052 <= 196059;
    i_distance_0053 <= 72414;
    i_distance_0054 <= 640098;
    i_distance_0055 <= 415717;
    i_distance_0056 <= 141547;
    i_distance_0057 <= 785389;
    i_distance_0058 <= 856305;
    i_distance_0059 <= 435829;
    i_distance_0060 <= 491381;
    i_distance_0061 <= 612343;
    i_distance_0062 <= 49659;
    i_distance_0063 <= 833535;
    correct_answer <= 9230;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 197764;
    i_distance_0001 <= 100485;
    i_distance_0002 <= 920582;
    i_distance_0003 <= 700935;
    i_distance_0004 <= 809352;
    i_distance_0005 <= 714758;
    i_distance_0006 <= 384138;
    i_distance_0007 <= 908556;
    i_distance_0008 <= 567053;
    i_distance_0009 <= 59022;
    i_distance_0010 <= 676370;
    i_distance_0011 <= 483986;
    i_distance_0012 <= 987156;
    i_distance_0013 <= 441111;
    i_distance_0014 <= 141080;
    i_distance_0015 <= 407833;
    i_distance_0016 <= 152473;
    i_distance_0017 <= 511133;
    i_distance_0018 <= 23198;
    i_distance_0019 <= 800507;
    i_distance_0020 <= 197152;
    i_distance_0021 <= 819105;
    i_distance_0022 <= 876834;
    i_distance_0023 <= 10148;
    i_distance_0024 <= 56741;
    i_distance_0025 <= 169895;
    i_distance_0026 <= 449581;
    i_distance_0027 <= 563763;
    i_distance_0028 <= 304565;
    i_distance_0029 <= 479031;
    i_distance_0030 <= 86456;
    i_distance_0031 <= 554039;
    i_distance_0032 <= 372027;
    i_distance_0033 <= 349506;
    i_distance_0034 <= 834242;
    i_distance_0035 <= 806340;
    i_distance_0036 <= 129734;
    i_distance_0037 <= 516678;
    i_distance_0038 <= 178378;
    i_distance_0039 <= 502859;
    i_distance_0040 <= 316106;
    i_distance_0041 <= 330317;
    i_distance_0042 <= 634186;
    i_distance_0043 <= 812106;
    i_distance_0044 <= 681041;
    i_distance_0045 <= 901717;
    i_distance_0046 <= 84310;
    i_distance_0047 <= 689750;
    i_distance_0048 <= 238040;
    i_distance_0049 <= 369880;
    i_distance_0050 <= 434269;
    i_distance_0051 <= 53345;
    i_distance_0052 <= 492517;
    i_distance_0053 <= 98151;
    i_distance_0054 <= 334697;
    i_distance_0055 <= 1025387;
    i_distance_0056 <= 785005;
    i_distance_0057 <= 967149;
    i_distance_0058 <= 510189;
    i_distance_0059 <= 27249;
    i_distance_0060 <= 71031;
    i_distance_0061 <= 78843;
    i_distance_0062 <= 1015037;
    i_distance_0063 <= 277118;
    correct_answer <= 10148;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 441219;
    i_distance_0001 <= 819973;
    i_distance_0002 <= 861829;
    i_distance_0003 <= 46983;
    i_distance_0004 <= 290693;
    i_distance_0005 <= 515335;
    i_distance_0006 <= 887814;
    i_distance_0007 <= 744587;
    i_distance_0008 <= 82699;
    i_distance_0009 <= 765199;
    i_distance_0010 <= 936080;
    i_distance_0011 <= 670866;
    i_distance_0012 <= 523411;
    i_distance_0013 <= 145433;
    i_distance_0014 <= 145434;
    i_distance_0015 <= 120473;
    i_distance_0016 <= 265758;
    i_distance_0017 <= 92831;
    i_distance_0018 <= 23842;
    i_distance_0019 <= 47010;
    i_distance_0020 <= 364196;
    i_distance_0021 <= 980262;
    i_distance_0022 <= 624168;
    i_distance_0023 <= 60459;
    i_distance_0024 <= 411436;
    i_distance_0025 <= 960047;
    i_distance_0026 <= 545584;
    i_distance_0027 <= 915508;
    i_distance_0028 <= 396982;
    i_distance_0029 <= 585530;
    i_distance_0030 <= 973115;
    i_distance_0031 <= 74171;
    i_distance_0032 <= 71229;
    i_distance_0033 <= 279230;
    i_distance_0034 <= 133694;
    i_distance_0035 <= 254912;
    i_distance_0036 <= 849091;
    i_distance_0037 <= 141895;
    i_distance_0038 <= 666448;
    i_distance_0039 <= 491605;
    i_distance_0040 <= 412630;
    i_distance_0041 <= 960471;
    i_distance_0042 <= 954197;
    i_distance_0043 <= 607324;
    i_distance_0044 <= 797922;
    i_distance_0045 <= 656483;
    i_distance_0046 <= 549478;
    i_distance_0047 <= 160103;
    i_distance_0048 <= 630505;
    i_distance_0049 <= 280170;
    i_distance_0050 <= 348906;
    i_distance_0051 <= 407018;
    i_distance_0052 <= 548333;
    i_distance_0053 <= 720878;
    i_distance_0054 <= 829678;
    i_distance_0055 <= 350187;
    i_distance_0056 <= 895474;
    i_distance_0057 <= 793588;
    i_distance_0058 <= 127477;
    i_distance_0059 <= 1040631;
    i_distance_0060 <= 696440;
    i_distance_0061 <= 1000442;
    i_distance_0062 <= 614908;
    i_distance_0063 <= 894589;
    correct_answer <= 23842;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 864641;
    i_distance_0001 <= 86529;
    i_distance_0002 <= 303234;
    i_distance_0003 <= 880516;
    i_distance_0004 <= 330629;
    i_distance_0005 <= 345095;
    i_distance_0006 <= 86154;
    i_distance_0007 <= 594065;
    i_distance_0008 <= 348434;
    i_distance_0009 <= 719893;
    i_distance_0010 <= 1011098;
    i_distance_0011 <= 875291;
    i_distance_0012 <= 874650;
    i_distance_0013 <= 828958;
    i_distance_0014 <= 345375;
    i_distance_0015 <= 826144;
    i_distance_0016 <= 628129;
    i_distance_0017 <= 716706;
    i_distance_0018 <= 773799;
    i_distance_0019 <= 70569;
    i_distance_0020 <= 851370;
    i_distance_0021 <= 993194;
    i_distance_0022 <= 35884;
    i_distance_0023 <= 1010733;
    i_distance_0024 <= 169898;
    i_distance_0025 <= 622767;
    i_distance_0026 <= 555953;
    i_distance_0027 <= 155703;
    i_distance_0028 <= 111544;
    i_distance_0029 <= 184505;
    i_distance_0030 <= 732092;
    i_distance_0031 <= 849724;
    i_distance_0032 <= 544190;
    i_distance_0033 <= 31807;
    i_distance_0034 <= 639804;
    i_distance_0035 <= 773825;
    i_distance_0036 <= 411076;
    i_distance_0037 <= 894148;
    i_distance_0038 <= 33861;
    i_distance_0039 <= 846788;
    i_distance_0040 <= 200393;
    i_distance_0041 <= 967882;
    i_distance_0042 <= 263243;
    i_distance_0043 <= 252627;
    i_distance_0044 <= 75988;
    i_distance_0045 <= 460887;
    i_distance_0046 <= 510935;
    i_distance_0047 <= 102105;
    i_distance_0048 <= 243034;
    i_distance_0049 <= 916186;
    i_distance_0050 <= 418017;
    i_distance_0051 <= 721252;
    i_distance_0052 <= 433764;
    i_distance_0053 <= 1007335;
    i_distance_0054 <= 248040;
    i_distance_0055 <= 879464;
    i_distance_0056 <= 97511;
    i_distance_0057 <= 972139;
    i_distance_0058 <= 834159;
    i_distance_0059 <= 496;
    i_distance_0060 <= 184819;
    i_distance_0061 <= 956916;
    i_distance_0062 <= 707701;
    i_distance_0063 <= 1028988;
    correct_answer <= 496;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 604289;
    i_distance_0001 <= 813186;
    i_distance_0002 <= 293123;
    i_distance_0003 <= 371202;
    i_distance_0004 <= 777090;
    i_distance_0005 <= 939785;
    i_distance_0006 <= 555275;
    i_distance_0007 <= 329359;
    i_distance_0008 <= 52241;
    i_distance_0009 <= 1045138;
    i_distance_0010 <= 3222;
    i_distance_0011 <= 682777;
    i_distance_0012 <= 383770;
    i_distance_0013 <= 900123;
    i_distance_0014 <= 647836;
    i_distance_0015 <= 817827;
    i_distance_0016 <= 585382;
    i_distance_0017 <= 124075;
    i_distance_0018 <= 782892;
    i_distance_0019 <= 1014574;
    i_distance_0020 <= 795185;
    i_distance_0021 <= 417074;
    i_distance_0022 <= 585395;
    i_distance_0023 <= 554164;
    i_distance_0024 <= 814135;
    i_distance_0025 <= 646456;
    i_distance_0026 <= 75704;
    i_distance_0027 <= 946106;
    i_distance_0028 <= 147898;
    i_distance_0029 <= 162749;
    i_distance_0030 <= 102590;
    i_distance_0031 <= 438079;
    i_distance_0032 <= 396993;
    i_distance_0033 <= 618561;
    i_distance_0034 <= 926787;
    i_distance_0035 <= 266308;
    i_distance_0036 <= 662597;
    i_distance_0037 <= 784326;
    i_distance_0038 <= 354249;
    i_distance_0039 <= 842573;
    i_distance_0040 <= 742221;
    i_distance_0041 <= 70095;
    i_distance_0042 <= 422609;
    i_distance_0043 <= 1016401;
    i_distance_0044 <= 277201;
    i_distance_0045 <= 523990;
    i_distance_0046 <= 721239;
    i_distance_0047 <= 143448;
    i_distance_0048 <= 978391;
    i_distance_0049 <= 708570;
    i_distance_0050 <= 125788;
    i_distance_0051 <= 912737;
    i_distance_0052 <= 878689;
    i_distance_0053 <= 110307;
    i_distance_0054 <= 177381;
    i_distance_0055 <= 892135;
    i_distance_0056 <= 894952;
    i_distance_0057 <= 940523;
    i_distance_0058 <= 374251;
    i_distance_0059 <= 683886;
    i_distance_0060 <= 168943;
    i_distance_0061 <= 903279;
    i_distance_0062 <= 548466;
    i_distance_0063 <= 858875;
    correct_answer <= 3222;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 605440;
    i_distance_0001 <= 201862;
    i_distance_0002 <= 1006473;
    i_distance_0003 <= 8331;
    i_distance_0004 <= 719116;
    i_distance_0005 <= 560141;
    i_distance_0006 <= 445965;
    i_distance_0007 <= 834447;
    i_distance_0008 <= 234767;
    i_distance_0009 <= 213905;
    i_distance_0010 <= 972187;
    i_distance_0011 <= 64412;
    i_distance_0012 <= 117409;
    i_distance_0013 <= 502949;
    i_distance_0014 <= 753831;
    i_distance_0015 <= 369960;
    i_distance_0016 <= 880042;
    i_distance_0017 <= 338862;
    i_distance_0018 <= 132735;
    i_distance_0019 <= 971439;
    i_distance_0020 <= 939566;
    i_distance_0021 <= 453042;
    i_distance_0022 <= 880435;
    i_distance_0023 <= 153906;
    i_distance_0024 <= 346934;
    i_distance_0025 <= 252091;
    i_distance_0026 <= 1042363;
    i_distance_0027 <= 379711;
    i_distance_0028 <= 939712;
    i_distance_0029 <= 501952;
    i_distance_0030 <= 926530;
    i_distance_0031 <= 248512;
    i_distance_0032 <= 163268;
    i_distance_0033 <= 180803;
    i_distance_0034 <= 620228;
    i_distance_0035 <= 710215;
    i_distance_0036 <= 746828;
    i_distance_0037 <= 188493;
    i_distance_0038 <= 461391;
    i_distance_0039 <= 883792;
    i_distance_0040 <= 403281;
    i_distance_0041 <= 2771;
    i_distance_0042 <= 221268;
    i_distance_0043 <= 306556;
    i_distance_0044 <= 121817;
    i_distance_0045 <= 759130;
    i_distance_0046 <= 1044059;
    i_distance_0047 <= 10457;
    i_distance_0048 <= 965853;
    i_distance_0049 <= 507998;
    i_distance_0050 <= 940380;
    i_distance_0051 <= 121948;
    i_distance_0052 <= 333026;
    i_distance_0053 <= 953572;
    i_distance_0054 <= 396261;
    i_distance_0055 <= 906090;
    i_distance_0056 <= 474987;
    i_distance_0057 <= 313323;
    i_distance_0058 <= 136430;
    i_distance_0059 <= 267638;
    i_distance_0060 <= 380278;
    i_distance_0061 <= 446076;
    i_distance_0062 <= 328318;
    i_distance_0063 <= 11647;
    correct_answer <= 2771;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 902531;
    i_distance_0001 <= 594566;
    i_distance_0002 <= 882824;
    i_distance_0003 <= 191242;
    i_distance_0004 <= 746763;
    i_distance_0005 <= 868364;
    i_distance_0006 <= 786574;
    i_distance_0007 <= 78226;
    i_distance_0008 <= 379542;
    i_distance_0009 <= 403478;
    i_distance_0010 <= 177689;
    i_distance_0011 <= 78873;
    i_distance_0012 <= 152093;
    i_distance_0013 <= 1036063;
    i_distance_0014 <= 13345;
    i_distance_0015 <= 48674;
    i_distance_0016 <= 996771;
    i_distance_0017 <= 613156;
    i_distance_0018 <= 223779;
    i_distance_0019 <= 796580;
    i_distance_0020 <= 758311;
    i_distance_0021 <= 982568;
    i_distance_0022 <= 637098;
    i_distance_0023 <= 930603;
    i_distance_0024 <= 857386;
    i_distance_0025 <= 911917;
    i_distance_0026 <= 113710;
    i_distance_0027 <= 572980;
    i_distance_0028 <= 861621;
    i_distance_0029 <= 761654;
    i_distance_0030 <= 1003064;
    i_distance_0031 <= 419385;
    i_distance_0032 <= 815802;
    i_distance_0033 <= 739771;
    i_distance_0034 <= 594112;
    i_distance_0035 <= 360643;
    i_distance_0036 <= 592067;
    i_distance_0037 <= 479685;
    i_distance_0038 <= 33606;
    i_distance_0039 <= 97095;
    i_distance_0040 <= 925517;
    i_distance_0041 <= 212178;
    i_distance_0042 <= 749144;
    i_distance_0043 <= 639324;
    i_distance_0044 <= 157277;
    i_distance_0045 <= 841695;
    i_distance_0046 <= 84193;
    i_distance_0047 <= 231650;
    i_distance_0048 <= 415201;
    i_distance_0049 <= 367588;
    i_distance_0050 <= 21605;
    i_distance_0051 <= 711270;
    i_distance_0052 <= 289125;
    i_distance_0053 <= 778477;
    i_distance_0054 <= 876909;
    i_distance_0055 <= 916463;
    i_distance_0056 <= 835055;
    i_distance_0057 <= 56815;
    i_distance_0058 <= 265587;
    i_distance_0059 <= 832755;
    i_distance_0060 <= 741621;
    i_distance_0061 <= 137591;
    i_distance_0062 <= 662909;
    i_distance_0063 <= 477694;
    correct_answer <= 13345;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 258307;
    i_distance_0001 <= 817795;
    i_distance_0002 <= 955779;
    i_distance_0003 <= 663558;
    i_distance_0004 <= 1031566;
    i_distance_0005 <= 512018;
    i_distance_0006 <= 210323;
    i_distance_0007 <= 861716;
    i_distance_0008 <= 580631;
    i_distance_0009 <= 157211;
    i_distance_0010 <= 275739;
    i_distance_0011 <= 787868;
    i_distance_0012 <= 327198;
    i_distance_0013 <= 644383;
    i_distance_0014 <= 23584;
    i_distance_0015 <= 748579;
    i_distance_0016 <= 91940;
    i_distance_0017 <= 315557;
    i_distance_0018 <= 473257;
    i_distance_0019 <= 890538;
    i_distance_0020 <= 996137;
    i_distance_0021 <= 468988;
    i_distance_0022 <= 540590;
    i_distance_0023 <= 427694;
    i_distance_0024 <= 1036208;
    i_distance_0025 <= 241072;
    i_distance_0026 <= 716979;
    i_distance_0027 <= 202166;
    i_distance_0028 <= 876344;
    i_distance_0029 <= 1001401;
    i_distance_0030 <= 74296;
    i_distance_0031 <= 152125;
    i_distance_0032 <= 176192;
    i_distance_0033 <= 295238;
    i_distance_0034 <= 524743;
    i_distance_0035 <= 330824;
    i_distance_0036 <= 553161;
    i_distance_0037 <= 196043;
    i_distance_0038 <= 819404;
    i_distance_0039 <= 74575;
    i_distance_0040 <= 684115;
    i_distance_0041 <= 838484;
    i_distance_0042 <= 484695;
    i_distance_0043 <= 123224;
    i_distance_0044 <= 913112;
    i_distance_0045 <= 679517;
    i_distance_0046 <= 501086;
    i_distance_0047 <= 237661;
    i_distance_0048 <= 842719;
    i_distance_0049 <= 601313;
    i_distance_0050 <= 349156;
    i_distance_0051 <= 593383;
    i_distance_0052 <= 497896;
    i_distance_0053 <= 951531;
    i_distance_0054 <= 653291;
    i_distance_0055 <= 226930;
    i_distance_0056 <= 130674;
    i_distance_0057 <= 406643;
    i_distance_0058 <= 392438;
    i_distance_0059 <= 364407;
    i_distance_0060 <= 387704;
    i_distance_0061 <= 757370;
    i_distance_0062 <= 410108;
    i_distance_0063 <= 642302;
    correct_answer <= 23584;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 909699;
    i_distance_0001 <= 356874;
    i_distance_0002 <= 603659;
    i_distance_0003 <= 301452;
    i_distance_0004 <= 1031821;
    i_distance_0005 <= 159628;
    i_distance_0006 <= 634123;
    i_distance_0007 <= 213904;
    i_distance_0008 <= 279697;
    i_distance_0009 <= 913041;
    i_distance_0010 <= 407060;
    i_distance_0011 <= 188438;
    i_distance_0012 <= 454678;
    i_distance_0013 <= 857753;
    i_distance_0014 <= 746906;
    i_distance_0015 <= 411768;
    i_distance_0016 <= 770209;
    i_distance_0017 <= 698018;
    i_distance_0018 <= 107683;
    i_distance_0019 <= 217380;
    i_distance_0020 <= 677285;
    i_distance_0021 <= 1022502;
    i_distance_0022 <= 328873;
    i_distance_0023 <= 39209;
    i_distance_0024 <= 625196;
    i_distance_0025 <= 115885;
    i_distance_0026 <= 25645;
    i_distance_0027 <= 391221;
    i_distance_0028 <= 458934;
    i_distance_0029 <= 377527;
    i_distance_0030 <= 880444;
    i_distance_0031 <= 391741;
    i_distance_0032 <= 11453;
    i_distance_0033 <= 151486;
    i_distance_0034 <= 964416;
    i_distance_0035 <= 51267;
    i_distance_0036 <= 60741;
    i_distance_0037 <= 464838;
    i_distance_0038 <= 494022;
    i_distance_0039 <= 501705;
    i_distance_0040 <= 723017;
    i_distance_0041 <= 523338;
    i_distance_0042 <= 1038154;
    i_distance_0043 <= 195920;
    i_distance_0044 <= 924368;
    i_distance_0045 <= 626388;
    i_distance_0046 <= 558167;
    i_distance_0047 <= 86747;
    i_distance_0048 <= 1042653;
    i_distance_0049 <= 593629;
    i_distance_0050 <= 765021;
    i_distance_0051 <= 280161;
    i_distance_0052 <= 185699;
    i_distance_0053 <= 407268;
    i_distance_0054 <= 964455;
    i_distance_0055 <= 734056;
    i_distance_0056 <= 497385;
    i_distance_0057 <= 673128;
    i_distance_0058 <= 74986;
    i_distance_0059 <= 659050;
    i_distance_0060 <= 89073;
    i_distance_0061 <= 1036146;
    i_distance_0062 <= 540277;
    i_distance_0063 <= 124152;
    correct_answer <= 11453;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 356864;
    i_distance_0001 <= 507137;
    i_distance_0002 <= 544773;
    i_distance_0003 <= 574988;
    i_distance_0004 <= 889228;
    i_distance_0005 <= 588812;
    i_distance_0006 <= 494095;
    i_distance_0007 <= 138894;
    i_distance_0008 <= 455824;
    i_distance_0009 <= 373906;
    i_distance_0010 <= 700181;
    i_distance_0011 <= 565274;
    i_distance_0012 <= 445339;
    i_distance_0013 <= 259997;
    i_distance_0014 <= 875934;
    i_distance_0015 <= 164637;
    i_distance_0016 <= 601125;
    i_distance_0017 <= 209704;
    i_distance_0018 <= 127020;
    i_distance_0019 <= 342832;
    i_distance_0020 <= 410289;
    i_distance_0021 <= 791989;
    i_distance_0022 <= 159415;
    i_distance_0023 <= 789303;
    i_distance_0024 <= 249657;
    i_distance_0025 <= 559673;
    i_distance_0026 <= 151867;
    i_distance_0027 <= 353335;
    i_distance_0028 <= 219325;
    i_distance_0029 <= 368446;
    i_distance_0030 <= 740031;
    i_distance_0031 <= 904894;
    i_distance_0032 <= 187579;
    i_distance_0033 <= 738373;
    i_distance_0034 <= 542535;
    i_distance_0035 <= 396231;
    i_distance_0036 <= 948169;
    i_distance_0037 <= 803275;
    i_distance_0038 <= 458323;
    i_distance_0039 <= 323540;
    i_distance_0040 <= 187221;
    i_distance_0041 <= 1018071;
    i_distance_0042 <= 81752;
    i_distance_0043 <= 595929;
    i_distance_0044 <= 819547;
    i_distance_0045 <= 367964;
    i_distance_0046 <= 726236;
    i_distance_0047 <= 696284;
    i_distance_0048 <= 1014626;
    i_distance_0049 <= 794468;
    i_distance_0050 <= 426469;
    i_distance_0051 <= 1011430;
    i_distance_0052 <= 623719;
    i_distance_0053 <= 836841;
    i_distance_0054 <= 467690;
    i_distance_0055 <= 985195;
    i_distance_0056 <= 205931;
    i_distance_0057 <= 936300;
    i_distance_0058 <= 744301;
    i_distance_0059 <= 563817;
    i_distance_0060 <= 450033;
    i_distance_0061 <= 480499;
    i_distance_0062 <= 474874;
    i_distance_0063 <= 559869;
    correct_answer <= 81752;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 59136;
    i_distance_0001 <= 596864;
    i_distance_0002 <= 228226;
    i_distance_0003 <= 977924;
    i_distance_0004 <= 110724;
    i_distance_0005 <= 313098;
    i_distance_0006 <= 475659;
    i_distance_0007 <= 110476;
    i_distance_0008 <= 45834;
    i_distance_0009 <= 700170;
    i_distance_0010 <= 139407;
    i_distance_0011 <= 98064;
    i_distance_0012 <= 1033106;
    i_distance_0013 <= 852245;
    i_distance_0014 <= 627989;
    i_distance_0015 <= 865046;
    i_distance_0016 <= 456725;
    i_distance_0017 <= 385945;
    i_distance_0018 <= 3868;
    i_distance_0019 <= 762526;
    i_distance_0020 <= 330142;
    i_distance_0021 <= 308638;
    i_distance_0022 <= 717348;
    i_distance_0023 <= 542501;
    i_distance_0024 <= 414886;
    i_distance_0025 <= 217383;
    i_distance_0026 <= 664234;
    i_distance_0027 <= 847531;
    i_distance_0028 <= 927403;
    i_distance_0029 <= 1046062;
    i_distance_0030 <= 295858;
    i_distance_0031 <= 833333;
    i_distance_0032 <= 596155;
    i_distance_0033 <= 970558;
    i_distance_0034 <= 160191;
    i_distance_0035 <= 350787;
    i_distance_0036 <= 1025988;
    i_distance_0037 <= 5574;
    i_distance_0038 <= 497096;
    i_distance_0039 <= 545482;
    i_distance_0040 <= 881100;
    i_distance_0041 <= 131149;
    i_distance_0042 <= 873423;
    i_distance_0043 <= 254288;
    i_distance_0044 <= 425424;
    i_distance_0045 <= 401108;
    i_distance_0046 <= 478805;
    i_distance_0047 <= 557274;
    i_distance_0048 <= 365660;
    i_distance_0049 <= 109022;
    i_distance_0050 <= 716767;
    i_distance_0051 <= 648932;
    i_distance_0052 <= 428775;
    i_distance_0053 <= 496872;
    i_distance_0054 <= 1038185;
    i_distance_0055 <= 774247;
    i_distance_0056 <= 950891;
    i_distance_0057 <= 675180;
    i_distance_0058 <= 661101;
    i_distance_0059 <= 473966;
    i_distance_0060 <= 627561;
    i_distance_0061 <= 6900;
    i_distance_0062 <= 851445;
    i_distance_0063 <= 665723;
    correct_answer <= 3868;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 972803;
    i_distance_0001 <= 3844;
    i_distance_0002 <= 481413;
    i_distance_0003 <= 709766;
    i_distance_0004 <= 378377;
    i_distance_0005 <= 628879;
    i_distance_0006 <= 900496;
    i_distance_0007 <= 461714;
    i_distance_0008 <= 930838;
    i_distance_0009 <= 647191;
    i_distance_0010 <= 1006235;
    i_distance_0011 <= 85020;
    i_distance_0012 <= 640027;
    i_distance_0013 <= 378656;
    i_distance_0014 <= 895392;
    i_distance_0015 <= 84898;
    i_distance_0016 <= 166179;
    i_distance_0017 <= 1026339;
    i_distance_0018 <= 590117;
    i_distance_0019 <= 790441;
    i_distance_0020 <= 449834;
    i_distance_0021 <= 206893;
    i_distance_0022 <= 165296;
    i_distance_0023 <= 803505;
    i_distance_0024 <= 458290;
    i_distance_0025 <= 255282;
    i_distance_0026 <= 833972;
    i_distance_0027 <= 783797;
    i_distance_0028 <= 780214;
    i_distance_0029 <= 122935;
    i_distance_0030 <= 225976;
    i_distance_0031 <= 95038;
    i_distance_0032 <= 243008;
    i_distance_0033 <= 495808;
    i_distance_0034 <= 228419;
    i_distance_0035 <= 345413;
    i_distance_0036 <= 85320;
    i_distance_0037 <= 982217;
    i_distance_0038 <= 149706;
    i_distance_0039 <= 797387;
    i_distance_0040 <= 599121;
    i_distance_0041 <= 189395;
    i_distance_0042 <= 1039700;
    i_distance_0043 <= 800212;
    i_distance_0044 <= 647385;
    i_distance_0045 <= 12508;
    i_distance_0046 <= 874204;
    i_distance_0047 <= 241657;
    i_distance_0048 <= 978658;
    i_distance_0049 <= 560867;
    i_distance_0050 <= 505443;
    i_distance_0051 <= 526178;
    i_distance_0052 <= 587494;
    i_distance_0053 <= 780139;
    i_distance_0054 <= 1036910;
    i_distance_0055 <= 216558;
    i_distance_0056 <= 645491;
    i_distance_0057 <= 638710;
    i_distance_0058 <= 798199;
    i_distance_0059 <= 870392;
    i_distance_0060 <= 651641;
    i_distance_0061 <= 338298;
    i_distance_0062 <= 891388;
    i_distance_0063 <= 173055;
    correct_answer <= 3844;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 476673;
    i_distance_0001 <= 69640;
    i_distance_0002 <= 888968;
    i_distance_0003 <= 826249;
    i_distance_0004 <= 951691;
    i_distance_0005 <= 876173;
    i_distance_0006 <= 934159;
    i_distance_0007 <= 88463;
    i_distance_0008 <= 117008;
    i_distance_0009 <= 520848;
    i_distance_0010 <= 458263;
    i_distance_0011 <= 836759;
    i_distance_0012 <= 248730;
    i_distance_0013 <= 554910;
    i_distance_0014 <= 376350;
    i_distance_0015 <= 982817;
    i_distance_0016 <= 854818;
    i_distance_0017 <= 395172;
    i_distance_0018 <= 126757;
    i_distance_0019 <= 1033893;
    i_distance_0020 <= 952743;
    i_distance_0021 <= 916648;
    i_distance_0022 <= 416681;
    i_distance_0023 <= 1027113;
    i_distance_0024 <= 646572;
    i_distance_0025 <= 215672;
    i_distance_0026 <= 694445;
    i_distance_0027 <= 578095;
    i_distance_0028 <= 282544;
    i_distance_0029 <= 634797;
    i_distance_0030 <= 263730;
    i_distance_0031 <= 669747;
    i_distance_0032 <= 632877;
    i_distance_0033 <= 102446;
    i_distance_0034 <= 695213;
    i_distance_0035 <= 946617;
    i_distance_0036 <= 731834;
    i_distance_0037 <= 959547;
    i_distance_0038 <= 862526;
    i_distance_0039 <= 1046719;
    i_distance_0040 <= 56388;
    i_distance_0041 <= 629705;
    i_distance_0042 <= 314057;
    i_distance_0043 <= 670033;
    i_distance_0044 <= 789458;
    i_distance_0045 <= 764372;
    i_distance_0046 <= 296024;
    i_distance_0047 <= 100573;
    i_distance_0048 <= 408544;
    i_distance_0049 <= 243811;
    i_distance_0050 <= 5995;
    i_distance_0051 <= 863852;
    i_distance_0052 <= 498795;
    i_distance_0053 <= 231019;
    i_distance_0054 <= 103279;
    i_distance_0055 <= 91632;
    i_distance_0056 <= 582265;
    i_distance_0057 <= 207472;
    i_distance_0058 <= 215155;
    i_distance_0059 <= 785392;
    i_distance_0060 <= 321014;
    i_distance_0061 <= 491254;
    i_distance_0062 <= 874872;
    i_distance_0063 <= 64761;
    correct_answer <= 5995;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 281601;
    i_distance_0001 <= 595714;
    i_distance_0002 <= 738051;
    i_distance_0003 <= 1028996;
    i_distance_0004 <= 855178;
    i_distance_0005 <= 612618;
    i_distance_0006 <= 315914;
    i_distance_0007 <= 231181;
    i_distance_0008 <= 183437;
    i_distance_0009 <= 588432;
    i_distance_0010 <= 439420;
    i_distance_0011 <= 363666;
    i_distance_0012 <= 25749;
    i_distance_0013 <= 573974;
    i_distance_0014 <= 369686;
    i_distance_0015 <= 404502;
    i_distance_0016 <= 922267;
    i_distance_0017 <= 889120;
    i_distance_0018 <= 433569;
    i_distance_0019 <= 715428;
    i_distance_0020 <= 642471;
    i_distance_0021 <= 376874;
    i_distance_0022 <= 1037482;
    i_distance_0023 <= 214573;
    i_distance_0024 <= 960302;
    i_distance_0025 <= 536494;
    i_distance_0026 <= 352175;
    i_distance_0027 <= 382001;
    i_distance_0028 <= 289459;
    i_distance_0029 <= 1020980;
    i_distance_0030 <= 244918;
    i_distance_0031 <= 975802;
    i_distance_0032 <= 992058;
    i_distance_0033 <= 160955;
    i_distance_0034 <= 467644;
    i_distance_0035 <= 912699;
    i_distance_0036 <= 116545;
    i_distance_0037 <= 444098;
    i_distance_0038 <= 1031746;
    i_distance_0039 <= 655042;
    i_distance_0040 <= 204098;
    i_distance_0041 <= 697413;
    i_distance_0042 <= 442054;
    i_distance_0043 <= 351433;
    i_distance_0044 <= 936778;
    i_distance_0045 <= 766923;
    i_distance_0046 <= 996809;
    i_distance_0047 <= 41427;
    i_distance_0048 <= 786771;
    i_distance_0049 <= 413655;
    i_distance_0050 <= 299480;
    i_distance_0051 <= 691169;
    i_distance_0052 <= 267622;
    i_distance_0053 <= 98791;
    i_distance_0054 <= 19689;
    i_distance_0055 <= 700142;
    i_distance_0056 <= 660084;
    i_distance_0057 <= 590966;
    i_distance_0058 <= 544503;
    i_distance_0059 <= 12280;
    i_distance_0060 <= 524541;
    i_distance_0061 <= 412667;
    i_distance_0062 <= 938364;
    i_distance_0063 <= 481661;
    correct_answer <= 12280;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 834821;
    i_distance_0001 <= 458246;
    i_distance_0002 <= 104071;
    i_distance_0003 <= 227461;
    i_distance_0004 <= 83462;
    i_distance_0005 <= 527238;
    i_distance_0006 <= 974347;
    i_distance_0007 <= 354827;
    i_distance_0008 <= 330256;
    i_distance_0009 <= 38417;
    i_distance_0010 <= 90770;
    i_distance_0011 <= 589075;
    i_distance_0012 <= 390676;
    i_distance_0013 <= 783637;
    i_distance_0014 <= 923157;
    i_distance_0015 <= 806288;
    i_distance_0016 <= 310804;
    i_distance_0017 <= 697497;
    i_distance_0018 <= 509085;
    i_distance_0019 <= 473759;
    i_distance_0020 <= 886688;
    i_distance_0021 <= 283808;
    i_distance_0022 <= 799138;
    i_distance_0023 <= 443045;
    i_distance_0024 <= 351399;
    i_distance_0025 <= 906279;
    i_distance_0026 <= 344617;
    i_distance_0027 <= 128044;
    i_distance_0028 <= 28461;
    i_distance_0029 <= 672431;
    i_distance_0030 <= 536882;
    i_distance_0031 <= 614194;
    i_distance_0032 <= 619444;
    i_distance_0033 <= 748341;
    i_distance_0034 <= 884150;
    i_distance_0035 <= 142267;
    i_distance_0036 <= 104892;
    i_distance_0037 <= 818750;
    i_distance_0038 <= 991679;
    i_distance_0039 <= 102596;
    i_distance_0040 <= 467269;
    i_distance_0041 <= 615109;
    i_distance_0042 <= 80458;
    i_distance_0043 <= 720974;
    i_distance_0044 <= 94799;
    i_distance_0045 <= 41040;
    i_distance_0046 <= 1041873;
    i_distance_0047 <= 978640;
    i_distance_0048 <= 763731;
    i_distance_0049 <= 468946;
    i_distance_0050 <= 1036886;
    i_distance_0051 <= 578396;
    i_distance_0052 <= 225887;
    i_distance_0053 <= 427106;
    i_distance_0054 <= 133603;
    i_distance_0055 <= 328293;
    i_distance_0056 <= 807662;
    i_distance_0057 <= 145520;
    i_distance_0058 <= 82291;
    i_distance_0059 <= 1036022;
    i_distance_0060 <= 13688;
    i_distance_0061 <= 355833;
    i_distance_0062 <= 237053;
    i_distance_0063 <= 836734;
    correct_answer <= 13688;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 1034880;
    i_distance_0001 <= 732678;
    i_distance_0002 <= 600329;
    i_distance_0003 <= 208394;
    i_distance_0004 <= 917386;
    i_distance_0005 <= 727180;
    i_distance_0006 <= 353041;
    i_distance_0007 <= 342674;
    i_distance_0008 <= 91545;
    i_distance_0009 <= 811808;
    i_distance_0010 <= 493861;
    i_distance_0011 <= 492198;
    i_distance_0012 <= 549544;
    i_distance_0013 <= 14248;
    i_distance_0014 <= 543791;
    i_distance_0015 <= 469167;
    i_distance_0016 <= 394161;
    i_distance_0017 <= 1033393;
    i_distance_0018 <= 466868;
    i_distance_0019 <= 457655;
    i_distance_0020 <= 824375;
    i_distance_0021 <= 619449;
    i_distance_0022 <= 461889;
    i_distance_0023 <= 238401;
    i_distance_0024 <= 48708;
    i_distance_0025 <= 965189;
    i_distance_0026 <= 731078;
    i_distance_0027 <= 658119;
    i_distance_0028 <= 167752;
    i_distance_0029 <= 856391;
    i_distance_0030 <= 875335;
    i_distance_0031 <= 48587;
    i_distance_0032 <= 289606;
    i_distance_0033 <= 369741;
    i_distance_0034 <= 764883;
    i_distance_0035 <= 813012;
    i_distance_0036 <= 253652;
    i_distance_0037 <= 934358;
    i_distance_0038 <= 262612;
    i_distance_0039 <= 8921;
    i_distance_0040 <= 578650;
    i_distance_0041 <= 1029851;
    i_distance_0042 <= 178140;
    i_distance_0043 <= 918748;
    i_distance_0044 <= 936935;
    i_distance_0045 <= 518121;
    i_distance_0046 <= 463594;
    i_distance_0047 <= 612971;
    i_distance_0048 <= 420460;
    i_distance_0049 <= 821997;
    i_distance_0050 <= 828654;
    i_distance_0051 <= 422767;
    i_distance_0052 <= 80753;
    i_distance_0053 <= 42354;
    i_distance_0054 <= 530164;
    i_distance_0055 <= 77813;
    i_distance_0056 <= 487157;
    i_distance_0057 <= 522871;
    i_distance_0058 <= 586489;
    i_distance_0059 <= 864634;
    i_distance_0060 <= 460283;
    i_distance_0061 <= 984829;
    i_distance_0062 <= 1024254;
    i_distance_0063 <= 169215;
    correct_answer <= 8921;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 968323;
    i_distance_0001 <= 1014277;
    i_distance_0002 <= 295558;
    i_distance_0003 <= 237447;
    i_distance_0004 <= 165241;
    i_distance_0005 <= 977674;
    i_distance_0006 <= 493324;
    i_distance_0007 <= 783887;
    i_distance_0008 <= 863889;
    i_distance_0009 <= 147346;
    i_distance_0010 <= 252307;
    i_distance_0011 <= 508692;
    i_distance_0012 <= 361877;
    i_distance_0013 <= 170134;
    i_distance_0014 <= 97047;
    i_distance_0015 <= 484630;
    i_distance_0016 <= 138136;
    i_distance_0017 <= 242586;
    i_distance_0018 <= 629144;
    i_distance_0019 <= 673686;
    i_distance_0020 <= 472989;
    i_distance_0021 <= 914974;
    i_distance_0022 <= 692001;
    i_distance_0023 <= 555044;
    i_distance_0024 <= 900389;
    i_distance_0025 <= 260773;
    i_distance_0026 <= 556330;
    i_distance_0027 <= 405549;
    i_distance_0028 <= 16816;
    i_distance_0029 <= 596528;
    i_distance_0030 <= 903088;
    i_distance_0031 <= 869300;
    i_distance_0032 <= 586549;
    i_distance_0033 <= 996151;
    i_distance_0034 <= 862903;
    i_distance_0035 <= 840248;
    i_distance_0036 <= 293432;
    i_distance_0037 <= 122816;
    i_distance_0038 <= 876355;
    i_distance_0039 <= 430275;
    i_distance_0040 <= 254024;
    i_distance_0041 <= 724427;
    i_distance_0042 <= 373835;
    i_distance_0043 <= 956755;
    i_distance_0044 <= 250069;
    i_distance_0045 <= 439765;
    i_distance_0046 <= 591703;
    i_distance_0047 <= 81403;
    i_distance_0048 <= 1006299;
    i_distance_0049 <= 170844;
    i_distance_0050 <= 709983;
    i_distance_0051 <= 838624;
    i_distance_0052 <= 549601;
    i_distance_0053 <= 616673;
    i_distance_0054 <= 874855;
    i_distance_0055 <= 600167;
    i_distance_0056 <= 140015;
    i_distance_0057 <= 122736;
    i_distance_0058 <= 58105;
    i_distance_0059 <= 349943;
    i_distance_0060 <= 598393;
    i_distance_0061 <= 1017595;
    i_distance_0062 <= 582141;
    i_distance_0063 <= 267134;
    correct_answer <= 16816;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 761858;
    i_distance_0001 <= 545539;
    i_distance_0002 <= 559363;
    i_distance_0003 <= 919049;
    i_distance_0004 <= 25481;
    i_distance_0005 <= 454929;
    i_distance_0006 <= 573972;
    i_distance_0007 <= 480789;
    i_distance_0008 <= 46998;
    i_distance_0009 <= 202903;
    i_distance_0010 <= 940948;
    i_distance_0011 <= 490772;
    i_distance_0012 <= 557082;
    i_distance_0013 <= 284188;
    i_distance_0014 <= 304285;
    i_distance_0015 <= 1032350;
    i_distance_0016 <= 109087;
    i_distance_0017 <= 988317;
    i_distance_0018 <= 13088;
    i_distance_0019 <= 43301;
    i_distance_0020 <= 949031;
    i_distance_0021 <= 502442;
    i_distance_0022 <= 773803;
    i_distance_0023 <= 489772;
    i_distance_0024 <= 399404;
    i_distance_0025 <= 426796;
    i_distance_0026 <= 380075;
    i_distance_0027 <= 769197;
    i_distance_0028 <= 614705;
    i_distance_0029 <= 992820;
    i_distance_0030 <= 1042740;
    i_distance_0031 <= 680502;
    i_distance_0032 <= 866744;
    i_distance_0033 <= 743609;
    i_distance_0034 <= 914233;
    i_distance_0035 <= 655803;
    i_distance_0036 <= 384316;
    i_distance_0037 <= 290237;
    i_distance_0038 <= 698172;
    i_distance_0039 <= 1042879;
    i_distance_0040 <= 914242;
    i_distance_0041 <= 15298;
    i_distance_0042 <= 853316;
    i_distance_0043 <= 347845;
    i_distance_0044 <= 483787;
    i_distance_0045 <= 548812;
    i_distance_0046 <= 580814;
    i_distance_0047 <= 835538;
    i_distance_0048 <= 179070;
    i_distance_0049 <= 318296;
    i_distance_0050 <= 948198;
    i_distance_0051 <= 238440;
    i_distance_0052 <= 673129;
    i_distance_0053 <= 446314;
    i_distance_0054 <= 316777;
    i_distance_0055 <= 474988;
    i_distance_0056 <= 578413;
    i_distance_0057 <= 16370;
    i_distance_0058 <= 269300;
    i_distance_0059 <= 571637;
    i_distance_0060 <= 677748;
    i_distance_0061 <= 449784;
    i_distance_0062 <= 971388;
    i_distance_0063 <= 977022;
    correct_answer <= 13088;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 573313;
    i_distance_0001 <= 478210;
    i_distance_0002 <= 562053;
    i_distance_0003 <= 893706;
    i_distance_0004 <= 1030797;
    i_distance_0005 <= 180494;
    i_distance_0006 <= 785553;
    i_distance_0007 <= 369042;
    i_distance_0008 <= 637457;
    i_distance_0009 <= 990612;
    i_distance_0010 <= 146076;
    i_distance_0011 <= 363038;
    i_distance_0012 <= 364320;
    i_distance_0013 <= 120865;
    i_distance_0014 <= 590497;
    i_distance_0015 <= 51619;
    i_distance_0016 <= 425508;
    i_distance_0017 <= 427645;
    i_distance_0018 <= 826538;
    i_distance_0019 <= 344107;
    i_distance_0020 <= 644011;
    i_distance_0021 <= 559917;
    i_distance_0022 <= 665516;
    i_distance_0023 <= 599343;
    i_distance_0024 <= 662959;
    i_distance_0025 <= 355507;
    i_distance_0026 <= 699833;
    i_distance_0027 <= 603582;
    i_distance_0028 <= 382272;
    i_distance_0029 <= 403777;
    i_distance_0030 <= 296130;
    i_distance_0031 <= 283842;
    i_distance_0032 <= 434249;
    i_distance_0033 <= 643529;
    i_distance_0034 <= 297547;
    i_distance_0035 <= 526027;
    i_distance_0036 <= 479824;
    i_distance_0037 <= 445010;
    i_distance_0038 <= 289109;
    i_distance_0039 <= 82776;
    i_distance_0040 <= 601178;
    i_distance_0041 <= 95579;
    i_distance_0042 <= 742108;
    i_distance_0043 <= 254940;
    i_distance_0044 <= 264285;
    i_distance_0045 <= 831453;
    i_distance_0046 <= 218204;
    i_distance_0047 <= 30171;
    i_distance_0048 <= 972771;
    i_distance_0049 <= 449764;
    i_distance_0050 <= 752741;
    i_distance_0051 <= 192232;
    i_distance_0052 <= 111849;
    i_distance_0053 <= 27497;
    i_distance_0054 <= 528747;
    i_distance_0055 <= 58861;
    i_distance_0056 <= 798960;
    i_distance_0057 <= 499312;
    i_distance_0058 <= 339315;
    i_distance_0059 <= 433653;
    i_distance_0060 <= 591480;
    i_distance_0061 <= 237945;
    i_distance_0062 <= 820092;
    i_distance_0063 <= 330237;
    correct_answer <= 27497;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 61056;
    i_distance_0001 <= 769665;
    i_distance_0002 <= 1015043;
    i_distance_0003 <= 884744;
    i_distance_0004 <= 281097;
    i_distance_0005 <= 1015947;
    i_distance_0006 <= 416141;
    i_distance_0007 <= 170768;
    i_distance_0008 <= 362385;
    i_distance_0009 <= 410130;
    i_distance_0010 <= 357394;
    i_distance_0011 <= 539413;
    i_distance_0012 <= 834453;
    i_distance_0013 <= 772507;
    i_distance_0014 <= 464670;
    i_distance_0015 <= 277408;
    i_distance_0016 <= 956664;
    i_distance_0017 <= 1014304;
    i_distance_0018 <= 58784;
    i_distance_0019 <= 776228;
    i_distance_0020 <= 158758;
    i_distance_0021 <= 577834;
    i_distance_0022 <= 554026;
    i_distance_0023 <= 681647;
    i_distance_0024 <= 247088;
    i_distance_0025 <= 933170;
    i_distance_0026 <= 365234;
    i_distance_0027 <= 175799;
    i_distance_0028 <= 809533;
    i_distance_0029 <= 778047;
    i_distance_0030 <= 116032;
    i_distance_0031 <= 661955;
    i_distance_0032 <= 218948;
    i_distance_0033 <= 757059;
    i_distance_0034 <= 697412;
    i_distance_0035 <= 309191;
    i_distance_0036 <= 919496;
    i_distance_0037 <= 176202;
    i_distance_0038 <= 678219;
    i_distance_0039 <= 950861;
    i_distance_0040 <= 813776;
    i_distance_0041 <= 769617;
    i_distance_0042 <= 623954;
    i_distance_0043 <= 626773;
    i_distance_0044 <= 373078;
    i_distance_0045 <= 211033;
    i_distance_0046 <= 323678;
    i_distance_0047 <= 336226;
    i_distance_0048 <= 487652;
    i_distance_0049 <= 344549;
    i_distance_0050 <= 483943;
    i_distance_0051 <= 516455;
    i_distance_0052 <= 720231;
    i_distance_0053 <= 214634;
    i_distance_0054 <= 382951;
    i_distance_0055 <= 863983;
    i_distance_0056 <= 508273;
    i_distance_0057 <= 367987;
    i_distance_0058 <= 624501;
    i_distance_0059 <= 888822;
    i_distance_0060 <= 944759;
    i_distance_0061 <= 228598;
    i_distance_0062 <= 528510;
    i_distance_0063 <= 522366;
    correct_answer <= 58784;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 409346;
    i_distance_0001 <= 497923;
    i_distance_0002 <= 241284;
    i_distance_0003 <= 767624;
    i_distance_0004 <= 353418;
    i_distance_0005 <= 220299;
    i_distance_0006 <= 749453;
    i_distance_0007 <= 94734;
    i_distance_0008 <= 778254;
    i_distance_0009 <= 844560;
    i_distance_0010 <= 401811;
    i_distance_0011 <= 1021980;
    i_distance_0012 <= 658205;
    i_distance_0013 <= 742689;
    i_distance_0014 <= 379810;
    i_distance_0015 <= 77475;
    i_distance_0016 <= 73252;
    i_distance_0017 <= 503461;
    i_distance_0018 <= 209830;
    i_distance_0019 <= 348583;
    i_distance_0020 <= 575015;
    i_distance_0021 <= 989098;
    i_distance_0022 <= 313259;
    i_distance_0023 <= 508972;
    i_distance_0024 <= 275116;
    i_distance_0025 <= 338478;
    i_distance_0026 <= 98479;
    i_distance_0027 <= 308781;
    i_distance_0028 <= 922286;
    i_distance_0029 <= 438451;
    i_distance_0030 <= 939445;
    i_distance_0031 <= 543030;
    i_distance_0032 <= 720568;
    i_distance_0033 <= 174521;
    i_distance_0034 <= 73020;
    i_distance_0035 <= 256704;
    i_distance_0036 <= 807618;
    i_distance_0037 <= 307654;
    i_distance_0038 <= 13894;
    i_distance_0039 <= 229576;
    i_distance_0040 <= 171081;
    i_distance_0041 <= 1003851;
    i_distance_0042 <= 471115;
    i_distance_0043 <= 745934;
    i_distance_0044 <= 78801;
    i_distance_0045 <= 563156;
    i_distance_0046 <= 418777;
    i_distance_0047 <= 141148;
    i_distance_0048 <= 31583;
    i_distance_0049 <= 252511;
    i_distance_0050 <= 421729;
    i_distance_0051 <= 479714;
    i_distance_0052 <= 995170;
    i_distance_0053 <= 421349;
    i_distance_0054 <= 141158;
    i_distance_0055 <= 580456;
    i_distance_0056 <= 662892;
    i_distance_0057 <= 683901;
    i_distance_0058 <= 357102;
    i_distance_0059 <= 134896;
    i_distance_0060 <= 227063;
    i_distance_0061 <= 500344;
    i_distance_0062 <= 553597;
    i_distance_0063 <= 780159;
    correct_answer <= 13894;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 720257;
    i_distance_0001 <= 1015684;
    i_distance_0002 <= 786826;
    i_distance_0003 <= 918286;
    i_distance_0004 <= 61205;
    i_distance_0005 <= 968856;
    i_distance_0006 <= 207642;
    i_distance_0007 <= 658587;
    i_distance_0008 <= 732188;
    i_distance_0009 <= 407328;
    i_distance_0010 <= 981793;
    i_distance_0011 <= 647202;
    i_distance_0012 <= 236835;
    i_distance_0013 <= 999972;
    i_distance_0014 <= 341284;
    i_distance_0015 <= 332968;
    i_distance_0016 <= 892586;
    i_distance_0017 <= 1002283;
    i_distance_0018 <= 337196;
    i_distance_0019 <= 442410;
    i_distance_0020 <= 563245;
    i_distance_0021 <= 368176;
    i_distance_0022 <= 487217;
    i_distance_0023 <= 368497;
    i_distance_0024 <= 859317;
    i_distance_0025 <= 206905;
    i_distance_0026 <= 240571;
    i_distance_0027 <= 935484;
    i_distance_0028 <= 525245;
    i_distance_0029 <= 559934;
    i_distance_0030 <= 614719;
    i_distance_0031 <= 559809;
    i_distance_0032 <= 435654;
    i_distance_0033 <= 607686;
    i_distance_0034 <= 893128;
    i_distance_0035 <= 901578;
    i_distance_0036 <= 710987;
    i_distance_0037 <= 408652;
    i_distance_0038 <= 206806;
    i_distance_0039 <= 816728;
    i_distance_0040 <= 704731;
    i_distance_0041 <= 929759;
    i_distance_0042 <= 184288;
    i_distance_0043 <= 110048;
    i_distance_0044 <= 464484;
    i_distance_0045 <= 267371;
    i_distance_0046 <= 932204;
    i_distance_0047 <= 913005;
    i_distance_0048 <= 441070;
    i_distance_0049 <= 300015;
    i_distance_0050 <= 872560;
    i_distance_0051 <= 649456;
    i_distance_0052 <= 217594;
    i_distance_0053 <= 241394;
    i_distance_0054 <= 286192;
    i_distance_0055 <= 762612;
    i_distance_0056 <= 910070;
    i_distance_0057 <= 947571;
    i_distance_0058 <= 413816;
    i_distance_0059 <= 1020016;
    i_distance_0060 <= 879866;
    i_distance_0061 <= 706811;
    i_distance_0062 <= 267004;
    i_distance_0063 <= 1033341;
    correct_answer <= 61205;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 212227;
    i_distance_0001 <= 551687;
    i_distance_0002 <= 12679;
    i_distance_0003 <= 120461;
    i_distance_0004 <= 1041680;
    i_distance_0005 <= 992656;
    i_distance_0006 <= 160402;
    i_distance_0007 <= 13717;
    i_distance_0008 <= 630422;
    i_distance_0009 <= 637975;
    i_distance_0010 <= 936598;
    i_distance_0011 <= 955673;
    i_distance_0012 <= 913690;
    i_distance_0013 <= 272155;
    i_distance_0014 <= 565531;
    i_distance_0015 <= 1027998;
    i_distance_0016 <= 365728;
    i_distance_0017 <= 417441;
    i_distance_0018 <= 895907;
    i_distance_0019 <= 715556;
    i_distance_0020 <= 159269;
    i_distance_0021 <= 521770;
    i_distance_0022 <= 624177;
    i_distance_0023 <= 901302;
    i_distance_0024 <= 926136;
    i_distance_0025 <= 332217;
    i_distance_0026 <= 620732;
    i_distance_0027 <= 153404;
    i_distance_0028 <= 155582;
    i_distance_0029 <= 669757;
    i_distance_0030 <= 451645;
    i_distance_0031 <= 454337;
    i_distance_0032 <= 716738;
    i_distance_0033 <= 197186;
    i_distance_0034 <= 125638;
    i_distance_0035 <= 863818;
    i_distance_0036 <= 896589;
    i_distance_0037 <= 426709;
    i_distance_0038 <= 152150;
    i_distance_0039 <= 531287;
    i_distance_0040 <= 681432;
    i_distance_0041 <= 167261;
    i_distance_0042 <= 251101;
    i_distance_0043 <= 389729;
    i_distance_0044 <= 921826;
    i_distance_0045 <= 879331;
    i_distance_0046 <= 443365;
    i_distance_0047 <= 685158;
    i_distance_0048 <= 1031015;
    i_distance_0049 <= 358760;
    i_distance_0050 <= 373990;
    i_distance_0051 <= 641002;
    i_distance_0052 <= 686955;
    i_distance_0053 <= 296299;
    i_distance_0054 <= 350318;
    i_distance_0055 <= 746482;
    i_distance_0056 <= 101491;
    i_distance_0057 <= 434551;
    i_distance_0058 <= 804088;
    i_distance_0059 <= 980089;
    i_distance_0060 <= 207354;
    i_distance_0061 <= 787708;
    i_distance_0062 <= 451709;
    i_distance_0063 <= 924414;
    correct_answer <= 12679;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 36358;
    i_distance_0001 <= 594185;
    i_distance_0002 <= 5770;
    i_distance_0003 <= 916234;
    i_distance_0004 <= 236684;
    i_distance_0005 <= 805646;
    i_distance_0006 <= 267282;
    i_distance_0007 <= 994839;
    i_distance_0008 <= 588441;
    i_distance_0009 <= 357532;
    i_distance_0010 <= 867613;
    i_distance_0011 <= 991011;
    i_distance_0012 <= 802852;
    i_distance_0013 <= 390949;
    i_distance_0014 <= 807594;
    i_distance_0015 <= 180396;
    i_distance_0016 <= 289843;
    i_distance_0017 <= 915251;
    i_distance_0018 <= 284797;
    i_distance_0019 <= 54707;
    i_distance_0020 <= 428344;
    i_distance_0021 <= 613561;
    i_distance_0022 <= 564156;
    i_distance_0023 <= 721341;
    i_distance_0024 <= 439613;
    i_distance_0025 <= 561599;
    i_distance_0026 <= 549692;
    i_distance_0027 <= 314617;
    i_distance_0028 <= 86089;
    i_distance_0029 <= 820043;
    i_distance_0030 <= 333004;
    i_distance_0031 <= 814795;
    i_distance_0032 <= 850510;
    i_distance_0033 <= 941390;
    i_distance_0034 <= 1046352;
    i_distance_0035 <= 937938;
    i_distance_0036 <= 309973;
    i_distance_0037 <= 721879;
    i_distance_0038 <= 257627;
    i_distance_0039 <= 968158;
    i_distance_0040 <= 707550;
    i_distance_0041 <= 251231;
    i_distance_0042 <= 358369;
    i_distance_0043 <= 505057;
    i_distance_0044 <= 914787;
    i_distance_0045 <= 1042020;
    i_distance_0046 <= 156008;
    i_distance_0047 <= 26729;
    i_distance_0048 <= 976488;
    i_distance_0049 <= 58603;
    i_distance_0050 <= 519912;
    i_distance_0051 <= 16232;
    i_distance_0052 <= 770413;
    i_distance_0053 <= 313839;
    i_distance_0054 <= 264560;
    i_distance_0055 <= 605297;
    i_distance_0056 <= 164210;
    i_distance_0057 <= 829169;
    i_distance_0058 <= 162805;
    i_distance_0059 <= 682486;
    i_distance_0060 <= 316279;
    i_distance_0061 <= 950390;
    i_distance_0062 <= 954745;
    i_distance_0063 <= 742781;
    correct_answer <= 5770;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 247298;
    i_distance_0001 <= 999554;
    i_distance_0002 <= 67717;
    i_distance_0003 <= 906117;
    i_distance_0004 <= 499591;
    i_distance_0005 <= 892805;
    i_distance_0006 <= 808458;
    i_distance_0007 <= 123787;
    i_distance_0008 <= 767630;
    i_distance_0009 <= 640145;
    i_distance_0010 <= 789394;
    i_distance_0011 <= 910355;
    i_distance_0012 <= 452243;
    i_distance_0013 <= 550037;
    i_distance_0014 <= 875929;
    i_distance_0015 <= 912409;
    i_distance_0016 <= 963867;
    i_distance_0017 <= 791581;
    i_distance_0018 <= 789282;
    i_distance_0019 <= 759330;
    i_distance_0020 <= 697719;
    i_distance_0021 <= 79867;
    i_distance_0022 <= 866215;
    i_distance_0023 <= 860712;
    i_distance_0024 <= 372907;
    i_distance_0025 <= 647212;
    i_distance_0026 <= 622509;
    i_distance_0027 <= 372526;
    i_distance_0028 <= 408240;
    i_distance_0029 <= 907060;
    i_distance_0030 <= 527412;
    i_distance_0031 <= 949815;
    i_distance_0032 <= 758840;
    i_distance_0033 <= 817594;
    i_distance_0034 <= 773563;
    i_distance_0035 <= 318779;
    i_distance_0036 <= 587708;
    i_distance_0037 <= 251580;
    i_distance_0038 <= 948543;
    i_distance_0039 <= 185920;
    i_distance_0040 <= 48191;
    i_distance_0041 <= 164420;
    i_distance_0042 <= 950860;
    i_distance_0043 <= 976591;
    i_distance_0044 <= 297552;
    i_distance_0045 <= 554199;
    i_distance_0046 <= 717787;
    i_distance_0047 <= 279389;
    i_distance_0048 <= 476510;
    i_distance_0049 <= 373343;
    i_distance_0050 <= 141537;
    i_distance_0051 <= 555623;
    i_distance_0052 <= 930920;
    i_distance_0053 <= 806526;
    i_distance_0054 <= 615402;
    i_distance_0055 <= 958829;
    i_distance_0056 <= 672494;
    i_distance_0057 <= 924911;
    i_distance_0058 <= 577011;
    i_distance_0059 <= 86517;
    i_distance_0060 <= 210935;
    i_distance_0061 <= 522235;
    i_distance_0062 <= 51710;
    i_distance_0063 <= 1001855;
    correct_answer <= 48191;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 104578;
    i_distance_0001 <= 682628;
    i_distance_0002 <= 344582;
    i_distance_0003 <= 980615;
    i_distance_0004 <= 21768;
    i_distance_0005 <= 662667;
    i_distance_0006 <= 495889;
    i_distance_0007 <= 687124;
    i_distance_0008 <= 1017365;
    i_distance_0009 <= 624279;
    i_distance_0010 <= 570906;
    i_distance_0011 <= 294427;
    i_distance_0012 <= 664737;
    i_distance_0013 <= 803110;
    i_distance_0014 <= 849319;
    i_distance_0015 <= 940200;
    i_distance_0016 <= 565932;
    i_distance_0017 <= 189998;
    i_distance_0018 <= 583854;
    i_distance_0019 <= 499377;
    i_distance_0020 <= 194746;
    i_distance_0021 <= 996924;
    i_distance_0022 <= 135103;
    i_distance_0023 <= 477376;
    i_distance_0024 <= 474305;
    i_distance_0025 <= 854592;
    i_distance_0026 <= 791107;
    i_distance_0027 <= 234436;
    i_distance_0028 <= 371141;
    i_distance_0029 <= 943178;
    i_distance_0030 <= 637899;
    i_distance_0031 <= 683596;
    i_distance_0032 <= 244171;
    i_distance_0033 <= 858959;
    i_distance_0034 <= 569937;
    i_distance_0035 <= 224722;
    i_distance_0036 <= 629075;
    i_distance_0037 <= 462548;
    i_distance_0038 <= 565716;
    i_distance_0039 <= 79576;
    i_distance_0040 <= 181850;
    i_distance_0041 <= 390362;
    i_distance_0042 <= 43357;
    i_distance_0043 <= 193886;
    i_distance_0044 <= 538718;
    i_distance_0045 <= 396638;
    i_distance_0046 <= 657121;
    i_distance_0047 <= 1023458;
    i_distance_0048 <= 950239;
    i_distance_0049 <= 192226;
    i_distance_0050 <= 909285;
    i_distance_0051 <= 1006952;
    i_distance_0052 <= 1046760;
    i_distance_0053 <= 763112;
    i_distance_0054 <= 538347;
    i_distance_0055 <= 997100;
    i_distance_0056 <= 617965;
    i_distance_0057 <= 212973;
    i_distance_0058 <= 272623;
    i_distance_0059 <= 441968;
    i_distance_0060 <= 1012719;
    i_distance_0061 <= 340458;
    i_distance_0062 <= 328698;
    i_distance_0063 <= 1044477;
    correct_answer <= 21768;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 415872;
    i_distance_0001 <= 674176;
    i_distance_0002 <= 73089;
    i_distance_0003 <= 674435;
    i_distance_0004 <= 62339;
    i_distance_0005 <= 535685;
    i_distance_0006 <= 8707;
    i_distance_0007 <= 201477;
    i_distance_0008 <= 94730;
    i_distance_0009 <= 778636;
    i_distance_0010 <= 426381;
    i_distance_0011 <= 112396;
    i_distance_0012 <= 45712;
    i_distance_0013 <= 34450;
    i_distance_0014 <= 913940;
    i_distance_0015 <= 218133;
    i_distance_0016 <= 930710;
    i_distance_0017 <= 731287;
    i_distance_0018 <= 677880;
    i_distance_0019 <= 774296;
    i_distance_0020 <= 854136;
    i_distance_0021 <= 304541;
    i_distance_0022 <= 757792;
    i_distance_0023 <= 532898;
    i_distance_0024 <= 724006;
    i_distance_0025 <= 191015;
    i_distance_0026 <= 1014824;
    i_distance_0027 <= 220841;
    i_distance_0028 <= 684330;
    i_distance_0029 <= 251433;
    i_distance_0030 <= 556972;
    i_distance_0031 <= 356518;
    i_distance_0032 <= 6321;
    i_distance_0033 <= 555315;
    i_distance_0034 <= 737337;
    i_distance_0035 <= 732858;
    i_distance_0036 <= 8123;
    i_distance_0037 <= 599878;
    i_distance_0038 <= 546248;
    i_distance_0039 <= 570442;
    i_distance_0040 <= 527229;
    i_distance_0041 <= 671694;
    i_distance_0042 <= 122836;
    i_distance_0043 <= 457943;
    i_distance_0044 <= 423896;
    i_distance_0045 <= 554967;
    i_distance_0046 <= 703834;
    i_distance_0047 <= 935383;
    i_distance_0048 <= 110172;
    i_distance_0049 <= 426457;
    i_distance_0050 <= 324574;
    i_distance_0051 <= 940128;
    i_distance_0052 <= 343778;
    i_distance_0053 <= 710245;
    i_distance_0054 <= 138214;
    i_distance_0055 <= 1015912;
    i_distance_0056 <= 671977;
    i_distance_0057 <= 708841;
    i_distance_0058 <= 687083;
    i_distance_0059 <= 642544;
    i_distance_0060 <= 698226;
    i_distance_0061 <= 765815;
    i_distance_0062 <= 408568;
    i_distance_0063 <= 798461;
    correct_answer <= 6321;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 410240;
    i_distance_0001 <= 122753;
    i_distance_0002 <= 689409;
    i_distance_0003 <= 20481;
    i_distance_0004 <= 188295;
    i_distance_0005 <= 391943;
    i_distance_0006 <= 918919;
    i_distance_0007 <= 727311;
    i_distance_0008 <= 1014929;
    i_distance_0009 <= 548625;
    i_distance_0010 <= 269336;
    i_distance_0011 <= 379033;
    i_distance_0012 <= 381339;
    i_distance_0013 <= 328732;
    i_distance_0014 <= 448667;
    i_distance_0015 <= 1037087;
    i_distance_0016 <= 548769;
    i_distance_0017 <= 442275;
    i_distance_0018 <= 936740;
    i_distance_0019 <= 864293;
    i_distance_0020 <= 561702;
    i_distance_0021 <= 481187;
    i_distance_0022 <= 593065;
    i_distance_0023 <= 36139;
    i_distance_0024 <= 1042731;
    i_distance_0025 <= 792494;
    i_distance_0026 <= 438959;
    i_distance_0027 <= 994990;
    i_distance_0028 <= 1041714;
    i_distance_0029 <= 110645;
    i_distance_0030 <= 96313;
    i_distance_0031 <= 693946;
    i_distance_0032 <= 755002;
    i_distance_0033 <= 194491;
    i_distance_0034 <= 198845;
    i_distance_0035 <= 225602;
    i_distance_0036 <= 729667;
    i_distance_0037 <= 218179;
    i_distance_0038 <= 772165;
    i_distance_0039 <= 981189;
    i_distance_0040 <= 438343;
    i_distance_0041 <= 758594;
    i_distance_0042 <= 996553;
    i_distance_0043 <= 523211;
    i_distance_0044 <= 324942;
    i_distance_0045 <= 763471;
    i_distance_0046 <= 140366;
    i_distance_0047 <= 170195;
    i_distance_0048 <= 696406;
    i_distance_0049 <= 337367;
    i_distance_0050 <= 210264;
    i_distance_0051 <= 599768;
    i_distance_0052 <= 608732;
    i_distance_0053 <= 762338;
    i_distance_0054 <= 617060;
    i_distance_0055 <= 56423;
    i_distance_0056 <= 485738;
    i_distance_0057 <= 943724;
    i_distance_0058 <= 252269;
    i_distance_0059 <= 537584;
    i_distance_0060 <= 765426;
    i_distance_0061 <= 466674;
    i_distance_0062 <= 712437;
    i_distance_0063 <= 677370;
    correct_answer <= 20481;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 939909;
    i_distance_0001 <= 989318;
    i_distance_0002 <= 481671;
    i_distance_0003 <= 810760;
    i_distance_0004 <= 799881;
    i_distance_0005 <= 390521;
    i_distance_0006 <= 702219;
    i_distance_0007 <= 225673;
    i_distance_0008 <= 387599;
    i_distance_0009 <= 383507;
    i_distance_0010 <= 968211;
    i_distance_0011 <= 836243;
    i_distance_0012 <= 917270;
    i_distance_0013 <= 113942;
    i_distance_0014 <= 30874;
    i_distance_0015 <= 437152;
    i_distance_0016 <= 26016;
    i_distance_0017 <= 630690;
    i_distance_0018 <= 621347;
    i_distance_0019 <= 167329;
    i_distance_0020 <= 260260;
    i_distance_0021 <= 899754;
    i_distance_0022 <= 280363;
    i_distance_0023 <= 145456;
    i_distance_0024 <= 944188;
    i_distance_0025 <= 92733;
    i_distance_0026 <= 20797;
    i_distance_0027 <= 535231;
    i_distance_0028 <= 498753;
    i_distance_0029 <= 230980;
    i_distance_0030 <= 138948;
    i_distance_0031 <= 395078;
    i_distance_0032 <= 589894;
    i_distance_0033 <= 759879;
    i_distance_0034 <= 863945;
    i_distance_0035 <= 483019;
    i_distance_0036 <= 789068;
    i_distance_0037 <= 18637;
    i_distance_0038 <= 733393;
    i_distance_0039 <= 830929;
    i_distance_0040 <= 601558;
    i_distance_0041 <= 314199;
    i_distance_0042 <= 647641;
    i_distance_0043 <= 396762;
    i_distance_0044 <= 278367;
    i_distance_0045 <= 198624;
    i_distance_0046 <= 942946;
    i_distance_0047 <= 39782;
    i_distance_0048 <= 883559;
    i_distance_0049 <= 228968;
    i_distance_0050 <= 543593;
    i_distance_0051 <= 1130;
    i_distance_0052 <= 120810;
    i_distance_0053 <= 810861;
    i_distance_0054 <= 726509;
    i_distance_0055 <= 575854;
    i_distance_0056 <= 669809;
    i_distance_0057 <= 527603;
    i_distance_0058 <= 372725;
    i_distance_0059 <= 507254;
    i_distance_0060 <= 523509;
    i_distance_0061 <= 599033;
    i_distance_0062 <= 479612;
    i_distance_0063 <= 840319;
    correct_answer <= 1130;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 513923;
    i_distance_0001 <= 47624;
    i_distance_0002 <= 5385;
    i_distance_0003 <= 982153;
    i_distance_0004 <= 220938;
    i_distance_0005 <= 142356;
    i_distance_0006 <= 590740;
    i_distance_0007 <= 269719;
    i_distance_0008 <= 210843;
    i_distance_0009 <= 440349;
    i_distance_0010 <= 161182;
    i_distance_0011 <= 680223;
    i_distance_0012 <= 925601;
    i_distance_0013 <= 924833;
    i_distance_0014 <= 495655;
    i_distance_0015 <= 746536;
    i_distance_0016 <= 990376;
    i_distance_0017 <= 325803;
    i_distance_0018 <= 799408;
    i_distance_0019 <= 659889;
    i_distance_0020 <= 221362;
    i_distance_0021 <= 357556;
    i_distance_0022 <= 686902;
    i_distance_0023 <= 407862;
    i_distance_0024 <= 27704;
    i_distance_0025 <= 977463;
    i_distance_0026 <= 9663;
    i_distance_0027 <= 1047743;
    i_distance_0028 <= 924225;
    i_distance_0029 <= 780994;
    i_distance_0030 <= 889535;
    i_distance_0031 <= 91716;
    i_distance_0032 <= 992581;
    i_distance_0033 <= 941515;
    i_distance_0034 <= 243022;
    i_distance_0035 <= 459343;
    i_distance_0036 <= 970193;
    i_distance_0037 <= 1006929;
    i_distance_0038 <= 520151;
    i_distance_0039 <= 417879;
    i_distance_0040 <= 180568;
    i_distance_0041 <= 299098;
    i_distance_0042 <= 81886;
    i_distance_0043 <= 886623;
    i_distance_0044 <= 408161;
    i_distance_0045 <= 1034722;
    i_distance_0046 <= 392295;
    i_distance_0047 <= 67305;
    i_distance_0048 <= 1036523;
    i_distance_0049 <= 341741;
    i_distance_0050 <= 634990;
    i_distance_0051 <= 368239;
    i_distance_0052 <= 827376;
    i_distance_0053 <= 24559;
    i_distance_0054 <= 510066;
    i_distance_0055 <= 489971;
    i_distance_0056 <= 163442;
    i_distance_0057 <= 549234;
    i_distance_0058 <= 634095;
    i_distance_0059 <= 879477;
    i_distance_0060 <= 955129;
    i_distance_0061 <= 413435;
    i_distance_0062 <= 644092;
    i_distance_0063 <= 126335;
    correct_answer <= 5385;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 701953;
    i_distance_0001 <= 395652;
    i_distance_0002 <= 174854;
    i_distance_0003 <= 786824;
    i_distance_0004 <= 86283;
    i_distance_0005 <= 737043;
    i_distance_0006 <= 148118;
    i_distance_0007 <= 497689;
    i_distance_0008 <= 18458;
    i_distance_0009 <= 160283;
    i_distance_0010 <= 83226;
    i_distance_0011 <= 891421;
    i_distance_0012 <= 583966;
    i_distance_0013 <= 395808;
    i_distance_0014 <= 557344;
    i_distance_0015 <= 414880;
    i_distance_0016 <= 388899;
    i_distance_0017 <= 530085;
    i_distance_0018 <= 571560;
    i_distance_0019 <= 813609;
    i_distance_0020 <= 844585;
    i_distance_0021 <= 25899;
    i_distance_0022 <= 1048109;
    i_distance_0023 <= 180528;
    i_distance_0024 <= 239153;
    i_distance_0025 <= 87728;
    i_distance_0026 <= 375989;
    i_distance_0027 <= 436662;
    i_distance_0028 <= 151864;
    i_distance_0029 <= 318136;
    i_distance_0030 <= 714682;
    i_distance_0031 <= 89788;
    i_distance_0032 <= 836797;
    i_distance_0033 <= 713534;
    i_distance_0034 <= 3134;
    i_distance_0035 <= 528065;
    i_distance_0036 <= 1039938;
    i_distance_0037 <= 341571;
    i_distance_0038 <= 256322;
    i_distance_0039 <= 269380;
    i_distance_0040 <= 703436;
    i_distance_0041 <= 885070;
    i_distance_0042 <= 863823;
    i_distance_0043 <= 88786;
    i_distance_0044 <= 86867;
    i_distance_0045 <= 238548;
    i_distance_0046 <= 1025108;
    i_distance_0047 <= 281302;
    i_distance_0048 <= 200919;
    i_distance_0049 <= 366809;
    i_distance_0050 <= 741337;
    i_distance_0051 <= 295132;
    i_distance_0052 <= 265189;
    i_distance_0053 <= 1024106;
    i_distance_0054 <= 306795;
    i_distance_0055 <= 547690;
    i_distance_0056 <= 755306;
    i_distance_0057 <= 766698;
    i_distance_0058 <= 180725;
    i_distance_0059 <= 236789;
    i_distance_0060 <= 551930;
    i_distance_0061 <= 187004;
    i_distance_0062 <= 577405;
    i_distance_0063 <= 8575;
    correct_answer <= 3134;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 164228;
    i_distance_0001 <= 131078;
    i_distance_0002 <= 227847;
    i_distance_0003 <= 167559;
    i_distance_0004 <= 96009;
    i_distance_0005 <= 540296;
    i_distance_0006 <= 258700;
    i_distance_0007 <= 1040269;
    i_distance_0008 <= 316174;
    i_distance_0009 <= 520078;
    i_distance_0010 <= 973712;
    i_distance_0011 <= 831376;
    i_distance_0012 <= 791182;
    i_distance_0013 <= 588428;
    i_distance_0014 <= 1008156;
    i_distance_0015 <= 59678;
    i_distance_0016 <= 917791;
    i_distance_0017 <= 732063;
    i_distance_0018 <= 242596;
    i_distance_0019 <= 734245;
    i_distance_0020 <= 325159;
    i_distance_0021 <= 1048104;
    i_distance_0022 <= 769712;
    i_distance_0023 <= 927280;
    i_distance_0024 <= 257072;
    i_distance_0025 <= 696242;
    i_distance_0026 <= 78900;
    i_distance_0027 <= 349365;
    i_distance_0028 <= 485430;
    i_distance_0029 <= 57399;
    i_distance_0030 <= 904375;
    i_distance_0031 <= 564407;
    i_distance_0032 <= 816442;
    i_distance_0033 <= 586172;
    i_distance_0034 <= 371648;
    i_distance_0035 <= 200768;
    i_distance_0036 <= 970946;
    i_distance_0037 <= 657477;
    i_distance_0038 <= 809597;
    i_distance_0039 <= 176198;
    i_distance_0040 <= 792269;
    i_distance_0041 <= 48591;
    i_distance_0042 <= 877396;
    i_distance_0043 <= 499925;
    i_distance_0044 <= 805208;
    i_distance_0045 <= 189018;
    i_distance_0046 <= 616796;
    i_distance_0047 <= 268895;
    i_distance_0048 <= 4836;
    i_distance_0049 <= 1024101;
    i_distance_0050 <= 217576;
    i_distance_0051 <= 501481;
    i_distance_0052 <= 609770;
    i_distance_0053 <= 545901;
    i_distance_0054 <= 648301;
    i_distance_0055 <= 415726;
    i_distance_0056 <= 128622;
    i_distance_0057 <= 282353;
    i_distance_0058 <= 782450;
    i_distance_0059 <= 127478;
    i_distance_0060 <= 271867;
    i_distance_0061 <= 1013629;
    i_distance_0062 <= 504574;
    i_distance_0063 <= 503167;
    correct_answer <= 4836;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 129536;
    i_distance_0001 <= 694532;
    i_distance_0002 <= 80772;
    i_distance_0003 <= 38788;
    i_distance_0004 <= 932235;
    i_distance_0005 <= 283276;
    i_distance_0006 <= 229007;
    i_distance_0007 <= 95635;
    i_distance_0008 <= 652948;
    i_distance_0009 <= 752533;
    i_distance_0010 <= 44565;
    i_distance_0011 <= 256409;
    i_distance_0012 <= 371738;
    i_distance_0013 <= 909594;
    i_distance_0014 <= 716697;
    i_distance_0015 <= 299161;
    i_distance_0016 <= 920094;
    i_distance_0017 <= 601881;
    i_distance_0018 <= 815903;
    i_distance_0019 <= 527009;
    i_distance_0020 <= 127648;
    i_distance_0021 <= 272421;
    i_distance_0022 <= 261419;
    i_distance_0023 <= 628779;
    i_distance_0024 <= 193580;
    i_distance_0025 <= 97711;
    i_distance_0026 <= 864562;
    i_distance_0027 <= 1005235;
    i_distance_0028 <= 566455;
    i_distance_0029 <= 156088;
    i_distance_0030 <= 717884;
    i_distance_0031 <= 539969;
    i_distance_0032 <= 219974;
    i_distance_0033 <= 61768;
    i_distance_0034 <= 651465;
    i_distance_0035 <= 202698;
    i_distance_0036 <= 792012;
    i_distance_0037 <= 881229;
    i_distance_0038 <= 136268;
    i_distance_0039 <= 733388;
    i_distance_0040 <= 550996;
    i_distance_0041 <= 629716;
    i_distance_0042 <= 186582;
    i_distance_0043 <= 666454;
    i_distance_0044 <= 216281;
    i_distance_0045 <= 162524;
    i_distance_0046 <= 809950;
    i_distance_0047 <= 114270;
    i_distance_0048 <= 506720;
    i_distance_0049 <= 375904;
    i_distance_0050 <= 285665;
    i_distance_0051 <= 949090;
    i_distance_0052 <= 1039844;
    i_distance_0053 <= 270331;
    i_distance_0054 <= 1020009;
    i_distance_0055 <= 730604;
    i_distance_0056 <= 215663;
    i_distance_0057 <= 781683;
    i_distance_0058 <= 525173;
    i_distance_0059 <= 795383;
    i_distance_0060 <= 213114;
    i_distance_0061 <= 960251;
    i_distance_0062 <= 585597;
    i_distance_0063 <= 364287;
    correct_answer <= 38788;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 40707;
    i_distance_0001 <= 634631;
    i_distance_0002 <= 235916;
    i_distance_0003 <= 809101;
    i_distance_0004 <= 315790;
    i_distance_0005 <= 810124;
    i_distance_0006 <= 699790;
    i_distance_0007 <= 627606;
    i_distance_0008 <= 408726;
    i_distance_0009 <= 160535;
    i_distance_0010 <= 511128;
    i_distance_0011 <= 997274;
    i_distance_0012 <= 977307;
    i_distance_0013 <= 608538;
    i_distance_0014 <= 392093;
    i_distance_0015 <= 806169;
    i_distance_0016 <= 159270;
    i_distance_0017 <= 8744;
    i_distance_0018 <= 538665;
    i_distance_0019 <= 226728;
    i_distance_0020 <= 261938;
    i_distance_0021 <= 606516;
    i_distance_0022 <= 370359;
    i_distance_0023 <= 778936;
    i_distance_0024 <= 251192;
    i_distance_0025 <= 24120;
    i_distance_0026 <= 526268;
    i_distance_0027 <= 758086;
    i_distance_0028 <= 979399;
    i_distance_0029 <= 992200;
    i_distance_0030 <= 349897;
    i_distance_0031 <= 367178;
    i_distance_0032 <= 330620;
    i_distance_0033 <= 973132;
    i_distance_0034 <= 917069;
    i_distance_0035 <= 293574;
    i_distance_0036 <= 206548;
    i_distance_0037 <= 466902;
    i_distance_0038 <= 745431;
    i_distance_0039 <= 95704;
    i_distance_0040 <= 733016;
    i_distance_0041 <= 229977;
    i_distance_0042 <= 470874;
    i_distance_0043 <= 84440;
    i_distance_0044 <= 352604;
    i_distance_0045 <= 526430;
    i_distance_0046 <= 713306;
    i_distance_0047 <= 665697;
    i_distance_0048 <= 1001187;
    i_distance_0049 <= 460259;
    i_distance_0050 <= 946789;
    i_distance_0051 <= 333414;
    i_distance_0052 <= 332903;
    i_distance_0053 <= 457447;
    i_distance_0054 <= 758889;
    i_distance_0055 <= 606569;
    i_distance_0056 <= 689005;
    i_distance_0057 <= 479598;
    i_distance_0058 <= 501871;
    i_distance_0059 <= 497263;
    i_distance_0060 <= 763380;
    i_distance_0061 <= 778102;
    i_distance_0062 <= 758396;
    i_distance_0063 <= 588798;
    correct_answer <= 8744;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 608897;
    i_distance_0001 <= 350593;
    i_distance_0002 <= 61569;
    i_distance_0003 <= 100738;
    i_distance_0004 <= 202632;
    i_distance_0005 <= 435337;
    i_distance_0006 <= 46223;
    i_distance_0007 <= 416144;
    i_distance_0008 <= 857361;
    i_distance_0009 <= 255634;
    i_distance_0010 <= 583035;
    i_distance_0011 <= 667921;
    i_distance_0012 <= 604950;
    i_distance_0013 <= 129435;
    i_distance_0014 <= 531868;
    i_distance_0015 <= 12061;
    i_distance_0016 <= 475167;
    i_distance_0017 <= 708385;
    i_distance_0018 <= 581410;
    i_distance_0019 <= 45860;
    i_distance_0020 <= 193829;
    i_distance_0021 <= 619818;
    i_distance_0022 <= 62123;
    i_distance_0023 <= 394797;
    i_distance_0024 <= 565038;
    i_distance_0025 <= 200752;
    i_distance_0026 <= 884659;
    i_distance_0027 <= 547124;
    i_distance_0028 <= 258868;
    i_distance_0029 <= 86840;
    i_distance_0030 <= 315449;
    i_distance_0031 <= 498109;
    i_distance_0032 <= 269758;
    i_distance_0033 <= 789699;
    i_distance_0034 <= 711620;
    i_distance_0035 <= 888391;
    i_distance_0036 <= 519880;
    i_distance_0037 <= 1044171;
    i_distance_0038 <= 75212;
    i_distance_0039 <= 238542;
    i_distance_0040 <= 408910;
    i_distance_0041 <= 521936;
    i_distance_0042 <= 95697;
    i_distance_0043 <= 248270;
    i_distance_0044 <= 68180;
    i_distance_0045 <= 4309;
    i_distance_0046 <= 308950;
    i_distance_0047 <= 830039;
    i_distance_0048 <= 761693;
    i_distance_0049 <= 382814;
    i_distance_0050 <= 1014493;
    i_distance_0051 <= 751586;
    i_distance_0052 <= 325987;
    i_distance_0053 <= 325605;
    i_distance_0054 <= 901477;
    i_distance_0055 <= 956135;
    i_distance_0056 <= 366957;
    i_distance_0057 <= 755053;
    i_distance_0058 <= 369009;
    i_distance_0059 <= 242419;
    i_distance_0060 <= 685942;
    i_distance_0061 <= 899447;
    i_distance_0062 <= 848632;
    i_distance_0063 <= 288891;
    correct_answer <= 4309;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 23681;
    i_distance_0001 <= 419970;
    i_distance_0002 <= 915201;
    i_distance_0003 <= 1020673;
    i_distance_0004 <= 473730;
    i_distance_0005 <= 58886;
    i_distance_0006 <= 770564;
    i_distance_0007 <= 75785;
    i_distance_0008 <= 321931;
    i_distance_0009 <= 341004;
    i_distance_0010 <= 1016460;
    i_distance_0011 <= 556046;
    i_distance_0012 <= 175631;
    i_distance_0013 <= 466061;
    i_distance_0014 <= 837264;
    i_distance_0015 <= 672786;
    i_distance_0016 <= 697235;
    i_distance_0017 <= 678548;
    i_distance_0018 <= 462476;
    i_distance_0019 <= 548886;
    i_distance_0020 <= 1012504;
    i_distance_0021 <= 477977;
    i_distance_0022 <= 231195;
    i_distance_0023 <= 266652;
    i_distance_0024 <= 288287;
    i_distance_0025 <= 606624;
    i_distance_0026 <= 494624;
    i_distance_0027 <= 339872;
    i_distance_0028 <= 541099;
    i_distance_0029 <= 347307;
    i_distance_0030 <= 495405;
    i_distance_0031 <= 984750;
    i_distance_0032 <= 569901;
    i_distance_0033 <= 503728;
    i_distance_0034 <= 828209;
    i_distance_0035 <= 312113;
    i_distance_0036 <= 598335;
    i_distance_0037 <= 893122;
    i_distance_0038 <= 997315;
    i_distance_0039 <= 2246;
    i_distance_0040 <= 941382;
    i_distance_0041 <= 125897;
    i_distance_0042 <= 971596;
    i_distance_0043 <= 980434;
    i_distance_0044 <= 368724;
    i_distance_0045 <= 506708;
    i_distance_0046 <= 118998;
    i_distance_0047 <= 244184;
    i_distance_0048 <= 1034458;
    i_distance_0049 <= 212443;
    i_distance_0050 <= 558173;
    i_distance_0051 <= 585309;
    i_distance_0052 <= 493280;
    i_distance_0053 <= 12386;
    i_distance_0054 <= 459366;
    i_distance_0055 <= 792936;
    i_distance_0056 <= 1003881;
    i_distance_0057 <= 36330;
    i_distance_0058 <= 969194;
    i_distance_0059 <= 746866;
    i_distance_0060 <= 1007219;
    i_distance_0061 <= 137333;
    i_distance_0062 <= 393851;
    i_distance_0063 <= 560765;
    correct_answer <= 2246;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 170624;
    i_distance_0001 <= 311553;
    i_distance_0002 <= 635266;
    i_distance_0003 <= 849540;
    i_distance_0004 <= 383748;
    i_distance_0005 <= 125446;
    i_distance_0006 <= 116487;
    i_distance_0007 <= 35208;
    i_distance_0008 <= 80650;
    i_distance_0009 <= 17931;
    i_distance_0010 <= 730124;
    i_distance_0011 <= 774027;
    i_distance_0012 <= 383756;
    i_distance_0013 <= 767886;
    i_distance_0014 <= 635408;
    i_distance_0015 <= 953619;
    i_distance_0016 <= 549782;
    i_distance_0017 <= 516503;
    i_distance_0018 <= 865560;
    i_distance_0019 <= 295958;
    i_distance_0020 <= 392858;
    i_distance_0021 <= 168985;
    i_distance_0022 <= 870429;
    i_distance_0023 <= 308765;
    i_distance_0024 <= 757279;
    i_distance_0025 <= 490018;
    i_distance_0026 <= 969122;
    i_distance_0027 <= 207908;
    i_distance_0028 <= 662694;
    i_distance_0029 <= 961196;
    i_distance_0030 <= 15154;
    i_distance_0031 <= 809522;
    i_distance_0032 <= 574521;
    i_distance_0033 <= 471099;
    i_distance_0034 <= 935357;
    i_distance_0035 <= 736832;
    i_distance_0036 <= 237891;
    i_distance_0037 <= 1032901;
    i_distance_0038 <= 623945;
    i_distance_0039 <= 230090;
    i_distance_0040 <= 737868;
    i_distance_0041 <= 851921;
    i_distance_0042 <= 394324;
    i_distance_0043 <= 308181;
    i_distance_0044 <= 1028182;
    i_distance_0045 <= 126550;
    i_distance_0046 <= 776277;
    i_distance_0047 <= 920447;
    i_distance_0048 <= 61019;
    i_distance_0049 <= 439515;
    i_distance_0050 <= 489308;
    i_distance_0051 <= 25566;
    i_distance_0052 <= 973662;
    i_distance_0053 <= 328160;
    i_distance_0054 <= 21987;
    i_distance_0055 <= 890339;
    i_distance_0056 <= 164713;
    i_distance_0057 <= 41577;
    i_distance_0058 <= 532073;
    i_distance_0059 <= 280181;
    i_distance_0060 <= 133110;
    i_distance_0061 <= 42745;
    i_distance_0062 <= 543483;
    i_distance_0063 <= 121855;
    correct_answer <= 15154;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 109568;
    i_distance_0001 <= 595970;
    i_distance_0002 <= 2694;
    i_distance_0003 <= 386311;
    i_distance_0004 <= 732936;
    i_distance_0005 <= 973963;
    i_distance_0006 <= 510604;
    i_distance_0007 <= 123404;
    i_distance_0008 <= 501900;
    i_distance_0009 <= 825743;
    i_distance_0010 <= 809103;
    i_distance_0011 <= 550926;
    i_distance_0012 <= 225944;
    i_distance_0013 <= 97560;
    i_distance_0014 <= 449051;
    i_distance_0015 <= 99836;
    i_distance_0016 <= 861595;
    i_distance_0017 <= 615840;
    i_distance_0018 <= 7200;
    i_distance_0019 <= 820899;
    i_distance_0020 <= 211751;
    i_distance_0021 <= 888361;
    i_distance_0022 <= 1042428;
    i_distance_0023 <= 472621;
    i_distance_0024 <= 809390;
    i_distance_0025 <= 604976;
    i_distance_0026 <= 385459;
    i_distance_0027 <= 775093;
    i_distance_0028 <= 852279;
    i_distance_0029 <= 396088;
    i_distance_0030 <= 1040571;
    i_distance_0031 <= 301117;
    i_distance_0032 <= 380223;
    i_distance_0033 <= 874179;
    i_distance_0034 <= 74182;
    i_distance_0035 <= 31309;
    i_distance_0036 <= 832336;
    i_distance_0037 <= 337105;
    i_distance_0038 <= 85200;
    i_distance_0039 <= 137682;
    i_distance_0040 <= 488020;
    i_distance_0041 <= 506069;
    i_distance_0042 <= 313939;
    i_distance_0043 <= 1005020;
    i_distance_0044 <= 90332;
    i_distance_0045 <= 440926;
    i_distance_0046 <= 17244;
    i_distance_0047 <= 449760;
    i_distance_0048 <= 219493;
    i_distance_0049 <= 172268;
    i_distance_0050 <= 467309;
    i_distance_0051 <= 29166;
    i_distance_0052 <= 1001967;
    i_distance_0053 <= 852207;
    i_distance_0054 <= 365938;
    i_distance_0055 <= 355316;
    i_distance_0056 <= 895733;
    i_distance_0057 <= 546293;
    i_distance_0058 <= 263157;
    i_distance_0059 <= 674036;
    i_distance_0060 <= 730233;
    i_distance_0061 <= 451324;
    i_distance_0062 <= 1047293;
    i_distance_0063 <= 536318;
    correct_answer <= 2694;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 398464;
    i_distance_0001 <= 919427;
    i_distance_0002 <= 605448;
    i_distance_0003 <= 400905;
    i_distance_0004 <= 953864;
    i_distance_0005 <= 176907;
    i_distance_0006 <= 211724;
    i_distance_0007 <= 445326;
    i_distance_0008 <= 99215;
    i_distance_0009 <= 276115;
    i_distance_0010 <= 276756;
    i_distance_0011 <= 825624;
    i_distance_0012 <= 99609;
    i_distance_0013 <= 456602;
    i_distance_0014 <= 774552;
    i_distance_0015 <= 438298;
    i_distance_0016 <= 32665;
    i_distance_0017 <= 123814;
    i_distance_0018 <= 762664;
    i_distance_0019 <= 193963;
    i_distance_0020 <= 661548;
    i_distance_0021 <= 639405;
    i_distance_0022 <= 518062;
    i_distance_0023 <= 159918;
    i_distance_0024 <= 34232;
    i_distance_0025 <= 415545;
    i_distance_0026 <= 782138;
    i_distance_0027 <= 384829;
    i_distance_0028 <= 315325;
    i_distance_0029 <= 722752;
    i_distance_0030 <= 239813;
    i_distance_0031 <= 952008;
    i_distance_0032 <= 964169;
    i_distance_0033 <= 982474;
    i_distance_0034 <= 698698;
    i_distance_0035 <= 116940;
    i_distance_0036 <= 513612;
    i_distance_0037 <= 639310;
    i_distance_0038 <= 195529;
    i_distance_0039 <= 178897;
    i_distance_0040 <= 498130;
    i_distance_0041 <= 64209;
    i_distance_0042 <= 419410;
    i_distance_0043 <= 404054;
    i_distance_0044 <= 596951;
    i_distance_0045 <= 107483;
    i_distance_0046 <= 260573;
    i_distance_0047 <= 985309;
    i_distance_0048 <= 804575;
    i_distance_0049 <= 187488;
    i_distance_0050 <= 537833;
    i_distance_0051 <= 195435;
    i_distance_0052 <= 649452;
    i_distance_0053 <= 202989;
    i_distance_0054 <= 530030;
    i_distance_0055 <= 101102;
    i_distance_0056 <= 119405;
    i_distance_0057 <= 691570;
    i_distance_0058 <= 719474;
    i_distance_0059 <= 118644;
    i_distance_0060 <= 332408;
    i_distance_0061 <= 162298;
    i_distance_0062 <= 547580;
    i_distance_0063 <= 29311;
    correct_answer <= 29311;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 108032;
    i_distance_0001 <= 173057;
    i_distance_0002 <= 955521;
    i_distance_0003 <= 982532;
    i_distance_0004 <= 398596;
    i_distance_0005 <= 327685;
    i_distance_0006 <= 796036;
    i_distance_0007 <= 388104;
    i_distance_0008 <= 480013;
    i_distance_0009 <= 142610;
    i_distance_0010 <= 987925;
    i_distance_0011 <= 890005;
    i_distance_0012 <= 855198;
    i_distance_0013 <= 72223;
    i_distance_0014 <= 134305;
    i_distance_0015 <= 749217;
    i_distance_0016 <= 159656;
    i_distance_0017 <= 233130;
    i_distance_0018 <= 706090;
    i_distance_0019 <= 459822;
    i_distance_0020 <= 905007;
    i_distance_0021 <= 550321;
    i_distance_0022 <= 824499;
    i_distance_0023 <= 763700;
    i_distance_0024 <= 1014580;
    i_distance_0025 <= 532021;
    i_distance_0026 <= 519863;
    i_distance_0027 <= 235827;
    i_distance_0028 <= 718649;
    i_distance_0029 <= 134713;
    i_distance_0030 <= 221369;
    i_distance_0031 <= 479421;
    i_distance_0032 <= 827967;
    i_distance_0033 <= 531903;
    i_distance_0034 <= 882112;
    i_distance_0035 <= 632387;
    i_distance_0036 <= 565059;
    i_distance_0037 <= 13253;
    i_distance_0038 <= 276805;
    i_distance_0039 <= 831815;
    i_distance_0040 <= 553285;
    i_distance_0041 <= 422983;
    i_distance_0042 <= 1013706;
    i_distance_0043 <= 133586;
    i_distance_0044 <= 598232;
    i_distance_0045 <= 1036376;
    i_distance_0046 <= 759516;
    i_distance_0047 <= 999646;
    i_distance_0048 <= 39134;
    i_distance_0049 <= 1012448;
    i_distance_0050 <= 835936;
    i_distance_0051 <= 560610;
    i_distance_0052 <= 181987;
    i_distance_0053 <= 869222;
    i_distance_0054 <= 690413;
    i_distance_0055 <= 254577;
    i_distance_0056 <= 227061;
    i_distance_0057 <= 82681;
    i_distance_0058 <= 239861;
    i_distance_0059 <= 740089;
    i_distance_0060 <= 1018618;
    i_distance_0061 <= 434939;
    i_distance_0062 <= 891900;
    i_distance_0063 <= 891773;
    correct_answer <= 13253;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 1023745;
    i_distance_0001 <= 236161;
    i_distance_0002 <= 683533;
    i_distance_0003 <= 639760;
    i_distance_0004 <= 103312;
    i_distance_0005 <= 363411;
    i_distance_0006 <= 866963;
    i_distance_0007 <= 234773;
    i_distance_0008 <= 110614;
    i_distance_0009 <= 562455;
    i_distance_0010 <= 141431;
    i_distance_0011 <= 991253;
    i_distance_0012 <= 736282;
    i_distance_0013 <= 768021;
    i_distance_0014 <= 533022;
    i_distance_0015 <= 822304;
    i_distance_0016 <= 568352;
    i_distance_0017 <= 721825;
    i_distance_0018 <= 863395;
    i_distance_0019 <= 910627;
    i_distance_0020 <= 486694;
    i_distance_0021 <= 923303;
    i_distance_0022 <= 760360;
    i_distance_0023 <= 454697;
    i_distance_0024 <= 864042;
    i_distance_0025 <= 553003;
    i_distance_0026 <= 811561;
    i_distance_0027 <= 706097;
    i_distance_0028 <= 477491;
    i_distance_0029 <= 107444;
    i_distance_0030 <= 795956;
    i_distance_0031 <= 704054;
    i_distance_0032 <= 171447;
    i_distance_0033 <= 843703;
    i_distance_0034 <= 782138;
    i_distance_0035 <= 291899;
    i_distance_0036 <= 343100;
    i_distance_0037 <= 141118;
    i_distance_0038 <= 490559;
    i_distance_0039 <= 9280;
    i_distance_0040 <= 352193;
    i_distance_0041 <= 91075;
    i_distance_0042 <= 515907;
    i_distance_0043 <= 382922;
    i_distance_0044 <= 11213;
    i_distance_0045 <= 439377;
    i_distance_0046 <= 831569;
    i_distance_0047 <= 791761;
    i_distance_0048 <= 715092;
    i_distance_0049 <= 812885;
    i_distance_0050 <= 500566;
    i_distance_0051 <= 203352;
    i_distance_0052 <= 780634;
    i_distance_0053 <= 563675;
    i_distance_0054 <= 859104;
    i_distance_0055 <= 306920;
    i_distance_0056 <= 529897;
    i_distance_0057 <= 437996;
    i_distance_0058 <= 940143;
    i_distance_0059 <= 153973;
    i_distance_0060 <= 783223;
    i_distance_0061 <= 38651;
    i_distance_0062 <= 883069;
    i_distance_0063 <= 820350;
    correct_answer <= 9280;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 698241;
    i_distance_0001 <= 58369;
    i_distance_0002 <= 268545;
    i_distance_0003 <= 544004;
    i_distance_0004 <= 922882;
    i_distance_0005 <= 372620;
    i_distance_0006 <= 321550;
    i_distance_0007 <= 792974;
    i_distance_0008 <= 714519;
    i_distance_0009 <= 202520;
    i_distance_0010 <= 1004061;
    i_distance_0011 <= 59936;
    i_distance_0012 <= 979617;
    i_distance_0013 <= 926245;
    i_distance_0014 <= 941479;
    i_distance_0015 <= 234922;
    i_distance_0016 <= 490925;
    i_distance_0017 <= 553646;
    i_distance_0018 <= 591792;
    i_distance_0019 <= 94514;
    i_distance_0020 <= 185781;
    i_distance_0021 <= 847542;
    i_distance_0022 <= 811959;
    i_distance_0023 <= 460600;
    i_distance_0024 <= 861497;
    i_distance_0025 <= 1006011;
    i_distance_0026 <= 625596;
    i_distance_0027 <= 129468;
    i_distance_0028 <= 832961;
    i_distance_0029 <= 72387;
    i_distance_0030 <= 779972;
    i_distance_0031 <= 517699;
    i_distance_0032 <= 638022;
    i_distance_0033 <= 510024;
    i_distance_0034 <= 657097;
    i_distance_0035 <= 192458;
    i_distance_0036 <= 1013836;
    i_distance_0037 <= 733006;
    i_distance_0038 <= 55119;
    i_distance_0039 <= 581968;
    i_distance_0040 <= 535503;
    i_distance_0041 <= 719316;
    i_distance_0042 <= 855892;
    i_distance_0043 <= 235606;
    i_distance_0044 <= 532827;
    i_distance_0045 <= 583519;
    i_distance_0046 <= 1025762;
    i_distance_0047 <= 438883;
    i_distance_0048 <= 785892;
    i_distance_0049 <= 272872;
    i_distance_0050 <= 948201;
    i_distance_0051 <= 71402;
    i_distance_0052 <= 700908;
    i_distance_0053 <= 320877;
    i_distance_0054 <= 490093;
    i_distance_0055 <= 943854;
    i_distance_0056 <= 887152;
    i_distance_0057 <= 94192;
    i_distance_0058 <= 396789;
    i_distance_0059 <= 520950;
    i_distance_0060 <= 658295;
    i_distance_0061 <= 1031289;
    i_distance_0062 <= 77565;
    i_distance_0063 <= 304767;
    correct_answer <= 55119;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 1031044;
    i_distance_0001 <= 598281;
    i_distance_0002 <= 641931;
    i_distance_0003 <= 679822;
    i_distance_0004 <= 528144;
    i_distance_0005 <= 832658;
    i_distance_0006 <= 967959;
    i_distance_0007 <= 778904;
    i_distance_0008 <= 978458;
    i_distance_0009 <= 296732;
    i_distance_0010 <= 43421;
    i_distance_0011 <= 88862;
    i_distance_0012 <= 125983;
    i_distance_0013 <= 1013534;
    i_distance_0014 <= 434465;
    i_distance_0015 <= 931618;
    i_distance_0016 <= 575011;
    i_distance_0017 <= 8357;
    i_distance_0018 <= 847400;
    i_distance_0019 <= 288552;
    i_distance_0020 <= 207914;
    i_distance_0021 <= 246608;
    i_distance_0022 <= 590382;
    i_distance_0023 <= 31797;
    i_distance_0024 <= 520636;
    i_distance_0025 <= 194237;
    i_distance_0026 <= 1001794;
    i_distance_0027 <= 560838;
    i_distance_0028 <= 190535;
    i_distance_0029 <= 243400;
    i_distance_0030 <= 426698;
    i_distance_0031 <= 545611;
    i_distance_0032 <= 1001676;
    i_distance_0033 <= 672077;
    i_distance_0034 <= 444623;
    i_distance_0035 <= 659536;
    i_distance_0036 <= 959568;
    i_distance_0037 <= 266578;
    i_distance_0038 <= 1005522;
    i_distance_0039 <= 384468;
    i_distance_0040 <= 686160;
    i_distance_0041 <= 839124;
    i_distance_0042 <= 409046;
    i_distance_0043 <= 793814;
    i_distance_0044 <= 859604;
    i_distance_0045 <= 291036;
    i_distance_0046 <= 605916;
    i_distance_0047 <= 783840;
    i_distance_0048 <= 120162;
    i_distance_0049 <= 738276;
    i_distance_0050 <= 377957;
    i_distance_0051 <= 234729;
    i_distance_0052 <= 335721;
    i_distance_0053 <= 980074;
    i_distance_0054 <= 409069;
    i_distance_0055 <= 272366;
    i_distance_0056 <= 913009;
    i_distance_0057 <= 408308;
    i_distance_0058 <= 455287;
    i_distance_0059 <= 941944;
    i_distance_0060 <= 867193;
    i_distance_0061 <= 658554;
    i_distance_0062 <= 143739;
    i_distance_0063 <= 570234;
    correct_answer <= 8357;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 919680;
    i_distance_0001 <= 257538;
    i_distance_0002 <= 33795;
    i_distance_0003 <= 872071;
    i_distance_0004 <= 675085;
    i_distance_0005 <= 862605;
    i_distance_0006 <= 267024;
    i_distance_0007 <= 615697;
    i_distance_0008 <= 266261;
    i_distance_0009 <= 459544;
    i_distance_0010 <= 513561;
    i_distance_0011 <= 377502;
    i_distance_0012 <= 231839;
    i_distance_0013 <= 261919;
    i_distance_0014 <= 547486;
    i_distance_0015 <= 760867;
    i_distance_0016 <= 428325;
    i_distance_0017 <= 801320;
    i_distance_0018 <= 698665;
    i_distance_0019 <= 608680;
    i_distance_0020 <= 878635;
    i_distance_0021 <= 702764;
    i_distance_0022 <= 727981;
    i_distance_0023 <= 977198;
    i_distance_0024 <= 157106;
    i_distance_0025 <= 38579;
    i_distance_0026 <= 201779;
    i_distance_0027 <= 232501;
    i_distance_0028 <= 781108;
    i_distance_0029 <= 883511;
    i_distance_0030 <= 403893;
    i_distance_0031 <= 795704;
    i_distance_0032 <= 187002;
    i_distance_0033 <= 1037885;
    i_distance_0034 <= 610878;
    i_distance_0035 <= 828992;
    i_distance_0036 <= 60481;
    i_distance_0037 <= 332226;
    i_distance_0038 <= 531396;
    i_distance_0039 <= 865220;
    i_distance_0040 <= 127559;
    i_distance_0041 <= 76999;
    i_distance_0042 <= 351100;
    i_distance_0043 <= 713291;
    i_distance_0044 <= 500556;
    i_distance_0045 <= 814541;
    i_distance_0046 <= 65617;
    i_distance_0047 <= 175828;
    i_distance_0048 <= 277846;
    i_distance_0049 <= 429054;
    i_distance_0050 <= 641881;
    i_distance_0051 <= 104667;
    i_distance_0052 <= 342236;
    i_distance_0053 <= 427485;
    i_distance_0054 <= 1044190;
    i_distance_0055 <= 141919;
    i_distance_0056 <= 45407;
    i_distance_0057 <= 549735;
    i_distance_0058 <= 1011191;
    i_distance_0059 <= 93560;
    i_distance_0060 <= 160378;
    i_distance_0061 <= 474235;
    i_distance_0062 <= 502524;
    i_distance_0063 <= 643966;
    correct_answer <= 33795;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 593024;
    i_distance_0001 <= 823808;
    i_distance_0002 <= 95107;
    i_distance_0003 <= 150404;
    i_distance_0004 <= 841989;
    i_distance_0005 <= 614281;
    i_distance_0006 <= 403726;
    i_distance_0007 <= 203919;
    i_distance_0008 <= 944526;
    i_distance_0009 <= 673274;
    i_distance_0010 <= 535955;
    i_distance_0011 <= 388118;
    i_distance_0012 <= 1038871;
    i_distance_0013 <= 77079;
    i_distance_0014 <= 518294;
    i_distance_0015 <= 448155;
    i_distance_0016 <= 847134;
    i_distance_0017 <= 963364;
    i_distance_0018 <= 576164;
    i_distance_0019 <= 726566;
    i_distance_0020 <= 355367;
    i_distance_0021 <= 616232;
    i_distance_0022 <= 864814;
    i_distance_0023 <= 658354;
    i_distance_0024 <= 595122;
    i_distance_0025 <= 960434;
    i_distance_0026 <= 252471;
    i_distance_0027 <= 51896;
    i_distance_0028 <= 677560;
    i_distance_0029 <= 708665;
    i_distance_0030 <= 198455;
    i_distance_0031 <= 288324;
    i_distance_0032 <= 122052;
    i_distance_0033 <= 1039046;
    i_distance_0034 <= 113353;
    i_distance_0035 <= 480201;
    i_distance_0036 <= 1000139;
    i_distance_0037 <= 100042;
    i_distance_0038 <= 453964;
    i_distance_0039 <= 756304;
    i_distance_0040 <= 80977;
    i_distance_0041 <= 619217;
    i_distance_0042 <= 522194;
    i_distance_0043 <= 998744;
    i_distance_0044 <= 793432;
    i_distance_0045 <= 198104;
    i_distance_0046 <= 295385;
    i_distance_0047 <= 995679;
    i_distance_0048 <= 678752;
    i_distance_0049 <= 710243;
    i_distance_0050 <= 517348;
    i_distance_0051 <= 980452;
    i_distance_0052 <= 530150;
    i_distance_0053 <= 603623;
    i_distance_0054 <= 498411;
    i_distance_0055 <= 554220;
    i_distance_0056 <= 450683;
    i_distance_0057 <= 710510;
    i_distance_0058 <= 776943;
    i_distance_0059 <= 792687;
    i_distance_0060 <= 361713;
    i_distance_0061 <= 781291;
    i_distance_0062 <= 719098;
    i_distance_0063 <= 975483;
    correct_answer <= 51896;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 1031426;
    i_distance_0001 <= 521475;
    i_distance_0002 <= 117764;
    i_distance_0003 <= 584582;
    i_distance_0004 <= 325513;
    i_distance_0005 <= 958474;
    i_distance_0006 <= 814731;
    i_distance_0007 <= 166926;
    i_distance_0008 <= 369807;
    i_distance_0009 <= 977422;
    i_distance_0010 <= 151058;
    i_distance_0011 <= 124953;
    i_distance_0012 <= 748827;
    i_distance_0013 <= 867867;
    i_distance_0014 <= 996765;
    i_distance_0015 <= 596763;
    i_distance_0016 <= 937247;
    i_distance_0017 <= 467999;
    i_distance_0018 <= 608417;
    i_distance_0019 <= 94371;
    i_distance_0020 <= 1004707;
    i_distance_0021 <= 8876;
    i_distance_0022 <= 211884;
    i_distance_0023 <= 228397;
    i_distance_0024 <= 527150;
    i_distance_0025 <= 609584;
    i_distance_0026 <= 837296;
    i_distance_0027 <= 641074;
    i_distance_0028 <= 672306;
    i_distance_0029 <= 617271;
    i_distance_0030 <= 1022651;
    i_distance_0031 <= 336700;
    i_distance_0032 <= 545472;
    i_distance_0033 <= 907330;
    i_distance_0034 <= 522310;
    i_distance_0035 <= 958407;
    i_distance_0036 <= 172236;
    i_distance_0037 <= 1869;
    i_distance_0038 <= 881741;
    i_distance_0039 <= 773713;
    i_distance_0040 <= 499795;
    i_distance_0041 <= 77524;
    i_distance_0042 <= 380884;
    i_distance_0043 <= 294870;
    i_distance_0044 <= 852825;
    i_distance_0045 <= 206170;
    i_distance_0046 <= 773082;
    i_distance_0047 <= 731738;
    i_distance_0048 <= 505822;
    i_distance_0049 <= 274659;
    i_distance_0050 <= 155242;
    i_distance_0051 <= 667882;
    i_distance_0052 <= 688620;
    i_distance_0053 <= 683116;
    i_distance_0054 <= 23277;
    i_distance_0055 <= 587498;
    i_distance_0056 <= 473455;
    i_distance_0057 <= 553713;
    i_distance_0058 <= 825713;
    i_distance_0059 <= 788209;
    i_distance_0060 <= 606201;
    i_distance_0061 <= 242170;
    i_distance_0062 <= 762108;
    i_distance_0063 <= 307709;
    correct_answer <= 1869;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 537866;
    i_distance_0001 <= 295180;
    i_distance_0002 <= 343183;
    i_distance_0003 <= 802834;
    i_distance_0004 <= 605588;
    i_distance_0005 <= 237718;
    i_distance_0006 <= 140695;
    i_distance_0007 <= 254358;
    i_distance_0008 <= 194462;
    i_distance_0009 <= 786718;
    i_distance_0010 <= 818336;
    i_distance_0011 <= 414112;
    i_distance_0012 <= 404642;
    i_distance_0013 <= 765987;
    i_distance_0014 <= 386980;
    i_distance_0015 <= 229925;
    i_distance_0016 <= 85542;
    i_distance_0017 <= 320676;
    i_distance_0018 <= 56360;
    i_distance_0019 <= 271912;
    i_distance_0020 <= 250921;
    i_distance_0021 <= 883752;
    i_distance_0022 <= 965549;
    i_distance_0023 <= 889006;
    i_distance_0024 <= 785453;
    i_distance_0025 <= 340656;
    i_distance_0026 <= 809649;
    i_distance_0027 <= 580275;
    i_distance_0028 <= 224948;
    i_distance_0029 <= 639285;
    i_distance_0030 <= 363443;
    i_distance_0031 <= 331448;
    i_distance_0032 <= 892866;
    i_distance_0033 <= 476997;
    i_distance_0034 <= 462790;
    i_distance_0035 <= 862279;
    i_distance_0036 <= 41544;
    i_distance_0037 <= 793033;
    i_distance_0038 <= 174155;
    i_distance_0039 <= 890062;
    i_distance_0040 <= 301391;
    i_distance_0041 <= 411087;
    i_distance_0042 <= 861009;
    i_distance_0043 <= 580946;
    i_distance_0044 <= 942675;
    i_distance_0045 <= 713812;
    i_distance_0046 <= 1004762;
    i_distance_0047 <= 681179;
    i_distance_0048 <= 474332;
    i_distance_0049 <= 747999;
    i_distance_0050 <= 799200;
    i_distance_0051 <= 1021540;
    i_distance_0052 <= 461925;
    i_distance_0053 <= 767590;
    i_distance_0054 <= 762854;
    i_distance_0055 <= 200171;
    i_distance_0056 <= 880111;
    i_distance_0057 <= 411505;
    i_distance_0058 <= 716787;
    i_distance_0059 <= 49141;
    i_distance_0060 <= 597878;
    i_distance_0061 <= 714743;
    i_distance_0062 <= 458360;
    i_distance_0063 <= 517500;
    correct_answer <= 41544;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 531457;
    i_distance_0001 <= 893316;
    i_distance_0002 <= 266244;
    i_distance_0003 <= 946052;
    i_distance_0004 <= 747784;
    i_distance_0005 <= 749705;
    i_distance_0006 <= 48392;
    i_distance_0007 <= 302091;
    i_distance_0008 <= 923922;
    i_distance_0009 <= 854290;
    i_distance_0010 <= 211476;
    i_distance_0011 <= 704022;
    i_distance_0012 <= 26137;
    i_distance_0013 <= 605597;
    i_distance_0014 <= 797087;
    i_distance_0015 <= 687781;
    i_distance_0016 <= 451114;
    i_distance_0017 <= 508715;
    i_distance_0018 <= 220588;
    i_distance_0019 <= 270254;
    i_distance_0020 <= 671663;
    i_distance_0021 <= 246704;
    i_distance_0022 <= 651695;
    i_distance_0023 <= 507058;
    i_distance_0024 <= 101683;
    i_distance_0025 <= 248368;
    i_distance_0026 <= 932280;
    i_distance_0027 <= 548795;
    i_distance_0028 <= 609084;
    i_distance_0029 <= 297278;
    i_distance_0030 <= 65729;
    i_distance_0031 <= 579777;
    i_distance_0032 <= 707137;
    i_distance_0033 <= 244037;
    i_distance_0034 <= 1022405;
    i_distance_0035 <= 12744;
    i_distance_0036 <= 642425;
    i_distance_0037 <= 730959;
    i_distance_0038 <= 133201;
    i_distance_0039 <= 624595;
    i_distance_0040 <= 844117;
    i_distance_0041 <= 350550;
    i_distance_0042 <= 1018969;
    i_distance_0043 <= 344154;
    i_distance_0044 <= 11995;
    i_distance_0045 <= 434011;
    i_distance_0046 <= 321885;
    i_distance_0047 <= 244574;
    i_distance_0048 <= 144865;
    i_distance_0049 <= 903651;
    i_distance_0050 <= 388581;
    i_distance_0051 <= 768486;
    i_distance_0052 <= 563430;
    i_distance_0053 <= 8040;
    i_distance_0054 <= 204775;
    i_distance_0055 <= 425325;
    i_distance_0056 <= 908783;
    i_distance_0057 <= 604914;
    i_distance_0058 <= 688883;
    i_distance_0059 <= 955894;
    i_distance_0060 <= 856313;
    i_distance_0061 <= 904059;
    i_distance_0062 <= 17534;
    i_distance_0063 <= 572159;
    correct_answer <= 8040;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 615040;
    i_distance_0001 <= 199427;
    i_distance_0002 <= 375045;
    i_distance_0003 <= 774021;
    i_distance_0004 <= 616055;
    i_distance_0005 <= 46600;
    i_distance_0006 <= 355462;
    i_distance_0007 <= 1048458;
    i_distance_0008 <= 701832;
    i_distance_0009 <= 664586;
    i_distance_0010 <= 187784;
    i_distance_0011 <= 104334;
    i_distance_0012 <= 753936;
    i_distance_0013 <= 3729;
    i_distance_0014 <= 736146;
    i_distance_0015 <= 22802;
    i_distance_0016 <= 273554;
    i_distance_0017 <= 916247;
    i_distance_0018 <= 407832;
    i_distance_0019 <= 655897;
    i_distance_0020 <= 141977;
    i_distance_0021 <= 953497;
    i_distance_0022 <= 160540;
    i_distance_0023 <= 538275;
    i_distance_0024 <= 682794;
    i_distance_0025 <= 523054;
    i_distance_0026 <= 958515;
    i_distance_0027 <= 602805;
    i_distance_0028 <= 607415;
    i_distance_0029 <= 996537;
    i_distance_0030 <= 176057;
    i_distance_0031 <= 561856;
    i_distance_0032 <= 135489;
    i_distance_0033 <= 1037762;
    i_distance_0034 <= 928452;
    i_distance_0035 <= 133959;
    i_distance_0036 <= 416718;
    i_distance_0037 <= 573647;
    i_distance_0038 <= 42704;
    i_distance_0039 <= 326734;
    i_distance_0040 <= 915026;
    i_distance_0041 <= 294994;
    i_distance_0042 <= 134612;
    i_distance_0043 <= 742485;
    i_distance_0044 <= 435407;
    i_distance_0045 <= 614359;
    i_distance_0046 <= 131163;
    i_distance_0047 <= 632546;
    i_distance_0048 <= 810595;
    i_distance_0049 <= 58466;
    i_distance_0050 <= 165223;
    i_distance_0051 <= 271337;
    i_distance_0052 <= 969578;
    i_distance_0053 <= 366058;
    i_distance_0054 <= 462319;
    i_distance_0055 <= 962672;
    i_distance_0056 <= 778735;
    i_distance_0057 <= 798578;
    i_distance_0058 <= 704500;
    i_distance_0059 <= 513525;
    i_distance_0060 <= 147447;
    i_distance_0061 <= 933370;
    i_distance_0062 <= 487163;
    i_distance_0063 <= 542461;
    correct_answer <= 3729;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 878209;
    i_distance_0001 <= 189315;
    i_distance_0002 <= 1033095;
    i_distance_0003 <= 458376;
    i_distance_0004 <= 1011464;
    i_distance_0005 <= 440202;
    i_distance_0006 <= 46859;
    i_distance_0007 <= 310286;
    i_distance_0008 <= 1009679;
    i_distance_0009 <= 891664;
    i_distance_0010 <= 6675;
    i_distance_0011 <= 495892;
    i_distance_0012 <= 224668;
    i_distance_0013 <= 261533;
    i_distance_0014 <= 591264;
    i_distance_0015 <= 669857;
    i_distance_0016 <= 275490;
    i_distance_0017 <= 878114;
    i_distance_0018 <= 960164;
    i_distance_0019 <= 988835;
    i_distance_0020 <= 932389;
    i_distance_0021 <= 835623;
    i_distance_0022 <= 845352;
    i_distance_0023 <= 924712;
    i_distance_0024 <= 495402;
    i_distance_0025 <= 701998;
    i_distance_0026 <= 1016121;
    i_distance_0027 <= 131513;
    i_distance_0028 <= 293563;
    i_distance_0029 <= 256188;
    i_distance_0030 <= 311357;
    i_distance_0031 <= 677566;
    i_distance_0032 <= 62015;
    i_distance_0033 <= 199613;
    i_distance_0034 <= 432068;
    i_distance_0035 <= 954053;
    i_distance_0036 <= 263367;
    i_distance_0037 <= 1025352;
    i_distance_0038 <= 295497;
    i_distance_0039 <= 64464;
    i_distance_0040 <= 979409;
    i_distance_0041 <= 645459;
    i_distance_0042 <= 1018198;
    i_distance_0043 <= 285143;
    i_distance_0044 <= 439638;
    i_distance_0045 <= 33241;
    i_distance_0046 <= 789850;
    i_distance_0047 <= 336093;
    i_distance_0048 <= 668895;
    i_distance_0049 <= 260705;
    i_distance_0050 <= 220258;
    i_distance_0051 <= 969443;
    i_distance_0052 <= 834791;
    i_distance_0053 <= 384616;
    i_distance_0054 <= 71020;
    i_distance_0055 <= 875117;
    i_distance_0056 <= 1011568;
    i_distance_0057 <= 981491;
    i_distance_0058 <= 208499;
    i_distance_0059 <= 561909;
    i_distance_0060 <= 1011705;
    i_distance_0061 <= 1023229;
    i_distance_0062 <= 873342;
    i_distance_0063 <= 483327;
    correct_answer <= 6675;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 398720;
    i_distance_0001 <= 617732;
    i_distance_0002 <= 7685;
    i_distance_0003 <= 181768;
    i_distance_0004 <= 418568;
    i_distance_0005 <= 816137;
    i_distance_0006 <= 490248;
    i_distance_0007 <= 155790;
    i_distance_0008 <= 167182;
    i_distance_0009 <= 777872;
    i_distance_0010 <= 686738;
    i_distance_0011 <= 99347;
    i_distance_0012 <= 1040916;
    i_distance_0013 <= 390936;
    i_distance_0014 <= 639129;
    i_distance_0015 <= 503324;
    i_distance_0016 <= 892835;
    i_distance_0017 <= 217639;
    i_distance_0018 <= 202023;
    i_distance_0019 <= 831529;
    i_distance_0020 <= 753705;
    i_distance_0021 <= 652459;
    i_distance_0022 <= 868268;
    i_distance_0023 <= 577584;
    i_distance_0024 <= 679857;
    i_distance_0025 <= 285360;
    i_distance_0026 <= 128435;
    i_distance_0027 <= 504120;
    i_distance_0028 <= 1011384;
    i_distance_0029 <= 238907;
    i_distance_0030 <= 457788;
    i_distance_0031 <= 869440;
    i_distance_0032 <= 529345;
    i_distance_0033 <= 683842;
    i_distance_0034 <= 378179;
    i_distance_0035 <= 219206;
    i_distance_0036 <= 705991;
    i_distance_0037 <= 313160;
    i_distance_0038 <= 905802;
    i_distance_0039 <= 1040715;
    i_distance_0040 <= 570830;
    i_distance_0041 <= 136270;
    i_distance_0042 <= 592978;
    i_distance_0043 <= 599634;
    i_distance_0044 <= 991709;
    i_distance_0045 <= 679133;
    i_distance_0046 <= 828127;
    i_distance_0047 <= 675297;
    i_distance_0048 <= 360161;
    i_distance_0049 <= 595681;
    i_distance_0050 <= 5857;
    i_distance_0051 <= 31080;
    i_distance_0052 <= 123242;
    i_distance_0053 <= 160618;
    i_distance_0054 <= 219627;
    i_distance_0055 <= 986477;
    i_distance_0056 <= 403435;
    i_distance_0057 <= 398963;
    i_distance_0058 <= 105334;
    i_distance_0059 <= 543352;
    i_distance_0060 <= 89593;
    i_distance_0061 <= 337658;
    i_distance_0062 <= 321915;
    i_distance_0063 <= 730620;
    correct_answer <= 5857;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 99584;
    i_distance_0001 <= 547713;
    i_distance_0002 <= 617858;
    i_distance_0003 <= 767880;
    i_distance_0004 <= 613000;
    i_distance_0005 <= 453647;
    i_distance_0006 <= 642448;
    i_distance_0007 <= 448916;
    i_distance_0008 <= 280084;
    i_distance_0009 <= 172565;
    i_distance_0010 <= 377880;
    i_distance_0011 <= 613661;
    i_distance_0012 <= 776868;
    i_distance_0013 <= 169343;
    i_distance_0014 <= 551593;
    i_distance_0015 <= 818734;
    i_distance_0016 <= 82864;
    i_distance_0017 <= 507826;
    i_distance_0018 <= 815540;
    i_distance_0019 <= 719925;
    i_distance_0020 <= 968246;
    i_distance_0021 <= 745014;
    i_distance_0022 <= 464952;
    i_distance_0023 <= 35253;
    i_distance_0024 <= 303162;
    i_distance_0025 <= 583990;
    i_distance_0026 <= 304317;
    i_distance_0027 <= 854590;
    i_distance_0028 <= 826047;
    i_distance_0029 <= 884160;
    i_distance_0030 <= 263744;
    i_distance_0031 <= 532290;
    i_distance_0032 <= 761791;
    i_distance_0033 <= 728516;
    i_distance_0034 <= 358725;
    i_distance_0035 <= 658630;
    i_distance_0036 <= 1038917;
    i_distance_0037 <= 547910;
    i_distance_0038 <= 732613;
    i_distance_0039 <= 499405;
    i_distance_0040 <= 892110;
    i_distance_0041 <= 47437;
    i_distance_0042 <= 170705;
    i_distance_0043 <= 553044;
    i_distance_0044 <= 396117;
    i_distance_0045 <= 35547;
    i_distance_0046 <= 143453;
    i_distance_0047 <= 954974;
    i_distance_0048 <= 145501;
    i_distance_0049 <= 1022051;
    i_distance_0050 <= 423782;
    i_distance_0051 <= 553830;
    i_distance_0052 <= 958696;
    i_distance_0053 <= 969449;
    i_distance_0054 <= 451432;
    i_distance_0055 <= 233578;
    i_distance_0056 <= 429168;
    i_distance_0057 <= 254204;
    i_distance_0058 <= 977781;
    i_distance_0059 <= 252277;
    i_distance_0060 <= 624758;
    i_distance_0061 <= 664699;
    i_distance_0062 <= 993020;
    i_distance_0063 <= 260863;
    correct_answer <= 35253;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 1003522;
    i_distance_0001 <= 248963;
    i_distance_0002 <= 121223;
    i_distance_0003 <= 67978;
    i_distance_0004 <= 143883;
    i_distance_0005 <= 2703;
    i_distance_0006 <= 43536;
    i_distance_0007 <= 931093;
    i_distance_0008 <= 388245;
    i_distance_0009 <= 168213;
    i_distance_0010 <= 195352;
    i_distance_0011 <= 71452;
    i_distance_0012 <= 163996;
    i_distance_0013 <= 302111;
    i_distance_0014 <= 471585;
    i_distance_0015 <= 56742;
    i_distance_0016 <= 924071;
    i_distance_0017 <= 729256;
    i_distance_0018 <= 892072;
    i_distance_0019 <= 978729;
    i_distance_0020 <= 111787;
    i_distance_0021 <= 652590;
    i_distance_0022 <= 534577;
    i_distance_0023 <= 593073;
    i_distance_0024 <= 818870;
    i_distance_0025 <= 649783;
    i_distance_0026 <= 173624;
    i_distance_0027 <= 779194;
    i_distance_0028 <= 553532;
    i_distance_0029 <= 310717;
    i_distance_0030 <= 121148;
    i_distance_0031 <= 953792;
    i_distance_0032 <= 195393;
    i_distance_0033 <= 616900;
    i_distance_0034 <= 286281;
    i_distance_0035 <= 20043;
    i_distance_0036 <= 32332;
    i_distance_0037 <= 718029;
    i_distance_0038 <= 870990;
    i_distance_0039 <= 357967;
    i_distance_0040 <= 510668;
    i_distance_0041 <= 794193;
    i_distance_0042 <= 527187;
    i_distance_0043 <= 677844;
    i_distance_0044 <= 699221;
    i_distance_0045 <= 419287;
    i_distance_0046 <= 31198;
    i_distance_0047 <= 179809;
    i_distance_0048 <= 307682;
    i_distance_0049 <= 1044707;
    i_distance_0050 <= 809700;
    i_distance_0051 <= 768225;
    i_distance_0052 <= 599270;
    i_distance_0053 <= 468459;
    i_distance_0054 <= 140524;
    i_distance_0055 <= 637549;
    i_distance_0056 <= 995054;
    i_distance_0057 <= 100973;
    i_distance_0058 <= 156529;
    i_distance_0059 <= 653298;
    i_distance_0060 <= 986482;
    i_distance_0061 <= 805237;
    i_distance_0062 <= 540028;
    i_distance_0063 <= 954366;
    correct_answer <= 2703;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 1034240;
    i_distance_0001 <= 546817;
    i_distance_0002 <= 960768;
    i_distance_0003 <= 332673;
    i_distance_0004 <= 268673;
    i_distance_0005 <= 662789;
    i_distance_0006 <= 498438;
    i_distance_0007 <= 857863;
    i_distance_0008 <= 647;
    i_distance_0009 <= 269705;
    i_distance_0010 <= 20746;
    i_distance_0011 <= 164361;
    i_distance_0012 <= 978700;
    i_distance_0013 <= 889221;
    i_distance_0014 <= 397445;
    i_distance_0015 <= 542991;
    i_distance_0016 <= 311188;
    i_distance_0017 <= 610068;
    i_distance_0018 <= 528917;
    i_distance_0019 <= 326551;
    i_distance_0020 <= 496409;
    i_distance_0021 <= 1001882;
    i_distance_0022 <= 735261;
    i_distance_0023 <= 548253;
    i_distance_0024 <= 139167;
    i_distance_0025 <= 567584;
    i_distance_0026 <= 974630;
    i_distance_0027 <= 421934;
    i_distance_0028 <= 750126;
    i_distance_0029 <= 656823;
    i_distance_0030 <= 145084;
    i_distance_0031 <= 409789;
    i_distance_0032 <= 888766;
    i_distance_0033 <= 157251;
    i_distance_0034 <= 187971;
    i_distance_0035 <= 805317;
    i_distance_0036 <= 580679;
    i_distance_0037 <= 199112;
    i_distance_0038 <= 20170;
    i_distance_0039 <= 167243;
    i_distance_0040 <= 589902;
    i_distance_0041 <= 751310;
    i_distance_0042 <= 590670;
    i_distance_0043 <= 951758;
    i_distance_0044 <= 973653;
    i_distance_0045 <= 465881;
    i_distance_0046 <= 729948;
    i_distance_0047 <= 478812;
    i_distance_0048 <= 133981;
    i_distance_0049 <= 797920;
    i_distance_0050 <= 893412;
    i_distance_0051 <= 362853;
    i_distance_0052 <= 550758;
    i_distance_0053 <= 139626;
    i_distance_0054 <= 182635;
    i_distance_0055 <= 894190;
    i_distance_0056 <= 663665;
    i_distance_0057 <= 559221;
    i_distance_0058 <= 1021686;
    i_distance_0059 <= 292728;
    i_distance_0060 <= 858619;
    i_distance_0061 <= 1010300;
    i_distance_0062 <= 772477;
    i_distance_0063 <= 541951;
    correct_answer <= 647;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 1031680;
    i_distance_0001 <= 412545;
    i_distance_0002 <= 649984;
    i_distance_0003 <= 629251;
    i_distance_0004 <= 208898;
    i_distance_0005 <= 856582;
    i_distance_0006 <= 101127;
    i_distance_0007 <= 739464;
    i_distance_0008 <= 937353;
    i_distance_0009 <= 197514;
    i_distance_0010 <= 294537;
    i_distance_0011 <= 796682;
    i_distance_0012 <= 343943;
    i_distance_0013 <= 711058;
    i_distance_0014 <= 960405;
    i_distance_0015 <= 382997;
    i_distance_0016 <= 43159;
    i_distance_0017 <= 368794;
    i_distance_0018 <= 163611;
    i_distance_0019 <= 138141;
    i_distance_0020 <= 781085;
    i_distance_0021 <= 97567;
    i_distance_0022 <= 106023;
    i_distance_0023 <= 102568;
    i_distance_0024 <= 392107;
    i_distance_0025 <= 509484;
    i_distance_0026 <= 361393;
    i_distance_0027 <= 1003314;
    i_distance_0028 <= 62389;
    i_distance_0029 <= 295605;
    i_distance_0030 <= 332342;
    i_distance_0031 <= 734136;
    i_distance_0032 <= 283962;
    i_distance_0033 <= 435772;
    i_distance_0034 <= 106045;
    i_distance_0035 <= 943169;
    i_distance_0036 <= 422853;
    i_distance_0037 <= 233285;
    i_distance_0038 <= 821193;
    i_distance_0039 <= 991179;
    i_distance_0040 <= 110156;
    i_distance_0041 <= 624460;
    i_distance_0042 <= 431310;
    i_distance_0043 <= 12626;
    i_distance_0044 <= 213459;
    i_distance_0045 <= 699227;
    i_distance_0046 <= 892380;
    i_distance_0047 <= 454238;
    i_distance_0048 <= 791903;
    i_distance_0049 <= 342753;
    i_distance_0050 <= 819426;
    i_distance_0051 <= 994786;
    i_distance_0052 <= 500196;
    i_distance_0053 <= 517864;
    i_distance_0054 <= 1030506;
    i_distance_0055 <= 45931;
    i_distance_0056 <= 660844;
    i_distance_0057 <= 709738;
    i_distance_0058 <= 793328;
    i_distance_0059 <= 922994;
    i_distance_0060 <= 705653;
    i_distance_0061 <= 882166;
    i_distance_0062 <= 827640;
    i_distance_0063 <= 216318;
    correct_answer <= 12626;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 507650;
    i_distance_0001 <= 678147;
    i_distance_0002 <= 954116;
    i_distance_0003 <= 708100;
    i_distance_0004 <= 462985;
    i_distance_0005 <= 711434;
    i_distance_0006 <= 407563;
    i_distance_0007 <= 290709;
    i_distance_0008 <= 986134;
    i_distance_0009 <= 367767;
    i_distance_0010 <= 526233;
    i_distance_0011 <= 672923;
    i_distance_0012 <= 902172;
    i_distance_0013 <= 183837;
    i_distance_0014 <= 516510;
    i_distance_0015 <= 683935;
    i_distance_0016 <= 614946;
    i_distance_0017 <= 932773;
    i_distance_0018 <= 429606;
    i_distance_0019 <= 517158;
    i_distance_0020 <= 536492;
    i_distance_0021 <= 840750;
    i_distance_0022 <= 450735;
    i_distance_0023 <= 37937;
    i_distance_0024 <= 927411;
    i_distance_0025 <= 865203;
    i_distance_0026 <= 646197;
    i_distance_0027 <= 806455;
    i_distance_0028 <= 855096;
    i_distance_0029 <= 554425;
    i_distance_0030 <= 567994;
    i_distance_0031 <= 643001;
    i_distance_0032 <= 468284;
    i_distance_0033 <= 145855;
    i_distance_0034 <= 993218;
    i_distance_0035 <= 43586;
    i_distance_0036 <= 354756;
    i_distance_0037 <= 865860;
    i_distance_0038 <= 18758;
    i_distance_0039 <= 457927;
    i_distance_0040 <= 994760;
    i_distance_0041 <= 996041;
    i_distance_0042 <= 113990;
    i_distance_0043 <= 50760;
    i_distance_0044 <= 765006;
    i_distance_0045 <= 204623;
    i_distance_0046 <= 287826;
    i_distance_0047 <= 1034195;
    i_distance_0048 <= 877524;
    i_distance_0049 <= 473684;
    i_distance_0050 <= 572503;
    i_distance_0051 <= 168411;
    i_distance_0052 <= 1039579;
    i_distance_0053 <= 229341;
    i_distance_0054 <= 531550;
    i_distance_0055 <= 605565;
    i_distance_0056 <= 851934;
    i_distance_0057 <= 320483;
    i_distance_0058 <= 148718;
    i_distance_0059 <= 592622;
    i_distance_0060 <= 893045;
    i_distance_0061 <= 133367;
    i_distance_0062 <= 800893;
    i_distance_0063 <= 562551;
    correct_answer <= 18758;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 450944;
    i_distance_0001 <= 404482;
    i_distance_0002 <= 299012;
    i_distance_0003 <= 220805;
    i_distance_0004 <= 900870;
    i_distance_0005 <= 540677;
    i_distance_0006 <= 542856;
    i_distance_0007 <= 289032;
    i_distance_0008 <= 605578;
    i_distance_0009 <= 11787;
    i_distance_0010 <= 115977;
    i_distance_0011 <= 829453;
    i_distance_0012 <= 464270;
    i_distance_0013 <= 419855;
    i_distance_0014 <= 828048;
    i_distance_0015 <= 913038;
    i_distance_0016 <= 130703;
    i_distance_0017 <= 675857;
    i_distance_0018 <= 1005978;
    i_distance_0019 <= 999194;
    i_distance_0020 <= 430240;
    i_distance_0021 <= 723361;
    i_distance_0022 <= 113569;
    i_distance_0023 <= 426019;
    i_distance_0024 <= 53413;
    i_distance_0025 <= 755962;
    i_distance_0026 <= 792110;
    i_distance_0027 <= 931118;
    i_distance_0028 <= 42672;
    i_distance_0029 <= 211258;
    i_distance_0030 <= 884283;
    i_distance_0031 <= 544443;
    i_distance_0032 <= 371902;
    i_distance_0033 <= 148927;
    i_distance_0034 <= 135486;
    i_distance_0035 <= 110400;
    i_distance_0036 <= 937155;
    i_distance_0037 <= 847684;
    i_distance_0038 <= 791491;
    i_distance_0039 <= 499908;
    i_distance_0040 <= 923593;
    i_distance_0041 <= 54729;
    i_distance_0042 <= 586834;
    i_distance_0043 <= 377684;
    i_distance_0044 <= 1005909;
    i_distance_0045 <= 348630;
    i_distance_0046 <= 601305;
    i_distance_0047 <= 101722;
    i_distance_0048 <= 596313;
    i_distance_0049 <= 54364;
    i_distance_0050 <= 475233;
    i_distance_0051 <= 367716;
    i_distance_0052 <= 678118;
    i_distance_0053 <= 436613;
    i_distance_0054 <= 20072;
    i_distance_0055 <= 643688;
    i_distance_0056 <= 617322;
    i_distance_0057 <= 122349;
    i_distance_0058 <= 439918;
    i_distance_0059 <= 562925;
    i_distance_0060 <= 711664;
    i_distance_0061 <= 607474;
    i_distance_0062 <= 264570;
    i_distance_0063 <= 674556;
    correct_answer <= 11787;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 581507;
    i_distance_0001 <= 955011;
    i_distance_0002 <= 868869;
    i_distance_0003 <= 70918;
    i_distance_0004 <= 254983;
    i_distance_0005 <= 414472;
    i_distance_0006 <= 546953;
    i_distance_0007 <= 406154;
    i_distance_0008 <= 866571;
    i_distance_0009 <= 757514;
    i_distance_0010 <= 543117;
    i_distance_0011 <= 489995;
    i_distance_0012 <= 660623;
    i_distance_0013 <= 216976;
    i_distance_0014 <= 242580;
    i_distance_0015 <= 234264;
    i_distance_0016 <= 324505;
    i_distance_0017 <= 936088;
    i_distance_0018 <= 871581;
    i_distance_0019 <= 994848;
    i_distance_0020 <= 298017;
    i_distance_0021 <= 260261;
    i_distance_0022 <= 730150;
    i_distance_0023 <= 185642;
    i_distance_0024 <= 15403;
    i_distance_0025 <= 424237;
    i_distance_0026 <= 814638;
    i_distance_0027 <= 724016;
    i_distance_0028 <= 246578;
    i_distance_0029 <= 442168;
    i_distance_0030 <= 54713;
    i_distance_0031 <= 48314;
    i_distance_0032 <= 852025;
    i_distance_0033 <= 262464;
    i_distance_0034 <= 613953;
    i_distance_0035 <= 963778;
    i_distance_0036 <= 282946;
    i_distance_0037 <= 505540;
    i_distance_0038 <= 1032905;
    i_distance_0039 <= 110921;
    i_distance_0040 <= 754130;
    i_distance_0041 <= 203731;
    i_distance_0042 <= 285395;
    i_distance_0043 <= 230613;
    i_distance_0044 <= 192854;
    i_distance_0045 <= 642901;
    i_distance_0046 <= 179029;
    i_distance_0047 <= 386394;
    i_distance_0048 <= 561372;
    i_distance_0049 <= 990304;
    i_distance_0050 <= 267233;
    i_distance_0051 <= 485865;
    i_distance_0052 <= 788843;
    i_distance_0053 <= 48363;
    i_distance_0054 <= 102891;
    i_distance_0055 <= 68843;
    i_distance_0056 <= 18286;
    i_distance_0057 <= 315628;
    i_distance_0058 <= 402803;
    i_distance_0059 <= 644980;
    i_distance_0060 <= 310261;
    i_distance_0061 <= 842739;
    i_distance_0062 <= 917112;
    i_distance_0063 <= 890747;
    correct_answer <= 15403;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 411904;
    i_distance_0001 <= 24067;
    i_distance_0002 <= 585476;
    i_distance_0003 <= 388873;
    i_distance_0004 <= 398985;
    i_distance_0005 <= 103947;
    i_distance_0006 <= 1006349;
    i_distance_0007 <= 507406;
    i_distance_0008 <= 89229;
    i_distance_0009 <= 406033;
    i_distance_0010 <= 912916;
    i_distance_0011 <= 416533;
    i_distance_0012 <= 887190;
    i_distance_0013 <= 688663;
    i_distance_0014 <= 490915;
    i_distance_0015 <= 125604;
    i_distance_0016 <= 435623;
    i_distance_0017 <= 199848;
    i_distance_0018 <= 834983;
    i_distance_0019 <= 1038890;
    i_distance_0020 <= 233004;
    i_distance_0021 <= 569645;
    i_distance_0022 <= 739579;
    i_distance_0023 <= 1035441;
    i_distance_0024 <= 943284;
    i_distance_0025 <= 324278;
    i_distance_0026 <= 947127;
    i_distance_0027 <= 864568;
    i_distance_0028 <= 653626;
    i_distance_0029 <= 314172;
    i_distance_0030 <= 776766;
    i_distance_0031 <= 594623;
    i_distance_0032 <= 888641;
    i_distance_0033 <= 798915;
    i_distance_0034 <= 118726;
    i_distance_0035 <= 542920;
    i_distance_0036 <= 554057;
    i_distance_0037 <= 40264;
    i_distance_0038 <= 325451;
    i_distance_0039 <= 824271;
    i_distance_0040 <= 32977;
    i_distance_0041 <= 492113;
    i_distance_0042 <= 925907;
    i_distance_0043 <= 482645;
    i_distance_0044 <= 87637;
    i_distance_0045 <= 760152;
    i_distance_0046 <= 893529;
    i_distance_0047 <= 590557;
    i_distance_0048 <= 367584;
    i_distance_0049 <= 237793;
    i_distance_0050 <= 385018;
    i_distance_0051 <= 300644;
    i_distance_0052 <= 489189;
    i_distance_0053 <= 936039;
    i_distance_0054 <= 982889;
    i_distance_0055 <= 491242;
    i_distance_0056 <= 733162;
    i_distance_0057 <= 668526;
    i_distance_0058 <= 403699;
    i_distance_0059 <= 142837;
    i_distance_0060 <= 832245;
    i_distance_0061 <= 412537;
    i_distance_0062 <= 639610;
    i_distance_0063 <= 1000187;
    correct_answer <= 24067;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 393730;
    i_distance_0001 <= 636802;
    i_distance_0002 <= 1030019;
    i_distance_0003 <= 263045;
    i_distance_0004 <= 146566;
    i_distance_0005 <= 777731;
    i_distance_0006 <= 704776;
    i_distance_0007 <= 968834;
    i_distance_0008 <= 74890;
    i_distance_0009 <= 436619;
    i_distance_0010 <= 884493;
    i_distance_0011 <= 315149;
    i_distance_0012 <= 963471;
    i_distance_0013 <= 995088;
    i_distance_0014 <= 652561;
    i_distance_0015 <= 158483;
    i_distance_0016 <= 353173;
    i_distance_0017 <= 908695;
    i_distance_0018 <= 919320;
    i_distance_0019 <= 881306;
    i_distance_0020 <= 924445;
    i_distance_0021 <= 247967;
    i_distance_0022 <= 488351;
    i_distance_0023 <= 560546;
    i_distance_0024 <= 873122;
    i_distance_0025 <= 464681;
    i_distance_0026 <= 985897;
    i_distance_0027 <= 651435;
    i_distance_0028 <= 1043627;
    i_distance_0029 <= 742958;
    i_distance_0030 <= 140335;
    i_distance_0031 <= 291252;
    i_distance_0032 <= 418869;
    i_distance_0033 <= 502965;
    i_distance_0034 <= 310837;
    i_distance_0035 <= 268088;
    i_distance_0036 <= 202299;
    i_distance_0037 <= 757439;
    i_distance_0038 <= 854080;
    i_distance_0039 <= 63870;
    i_distance_0040 <= 684739;
    i_distance_0041 <= 413386;
    i_distance_0042 <= 278477;
    i_distance_0043 <= 867149;
    i_distance_0044 <= 704596;
    i_distance_0045 <= 976986;
    i_distance_0046 <= 1016030;
    i_distance_0047 <= 637919;
    i_distance_0048 <= 647010;
    i_distance_0049 <= 776035;
    i_distance_0050 <= 530534;
    i_distance_0051 <= 445160;
    i_distance_0052 <= 617837;
    i_distance_0053 <= 884590;
    i_distance_0054 <= 293103;
    i_distance_0055 <= 968688;
    i_distance_0056 <= 756461;
    i_distance_0057 <= 114035;
    i_distance_0058 <= 763380;
    i_distance_0059 <= 461815;
    i_distance_0060 <= 378873;
    i_distance_0061 <= 361083;
    i_distance_0062 <= 928892;
    i_distance_0063 <= 339582;
    correct_answer <= 63870;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 893313;
    i_distance_0001 <= 18818;
    i_distance_0002 <= 739843;
    i_distance_0003 <= 1041028;
    i_distance_0004 <= 226438;
    i_distance_0005 <= 316551;
    i_distance_0006 <= 15884;
    i_distance_0007 <= 1046797;
    i_distance_0008 <= 246286;
    i_distance_0009 <= 546830;
    i_distance_0010 <= 483984;
    i_distance_0011 <= 390412;
    i_distance_0012 <= 925200;
    i_distance_0013 <= 364691;
    i_distance_0014 <= 422807;
    i_distance_0015 <= 907799;
    i_distance_0016 <= 272793;
    i_distance_0017 <= 346008;
    i_distance_0018 <= 26908;
    i_distance_0019 <= 1013535;
    i_distance_0020 <= 307744;
    i_distance_0021 <= 908964;
    i_distance_0022 <= 55078;
    i_distance_0023 <= 205094;
    i_distance_0024 <= 981551;
    i_distance_0025 <= 220592;
    i_distance_0026 <= 671026;
    i_distance_0027 <= 247475;
    i_distance_0028 <= 608820;
    i_distance_0029 <= 963131;
    i_distance_0030 <= 183484;
    i_distance_0031 <= 390590;
    i_distance_0032 <= 467140;
    i_distance_0033 <= 58054;
    i_distance_0034 <= 482887;
    i_distance_0035 <= 207691;
    i_distance_0036 <= 934859;
    i_distance_0037 <= 905805;
    i_distance_0038 <= 975951;
    i_distance_0039 <= 449360;
    i_distance_0040 <= 427088;
    i_distance_0041 <= 415439;
    i_distance_0042 <= 834898;
    i_distance_0043 <= 595669;
    i_distance_0044 <= 433913;
    i_distance_0045 <= 201559;
    i_distance_0046 <= 526935;
    i_distance_0047 <= 477535;
    i_distance_0048 <= 398434;
    i_distance_0049 <= 719848;
    i_distance_0050 <= 770539;
    i_distance_0051 <= 813294;
    i_distance_0052 <= 281840;
    i_distance_0053 <= 355569;
    i_distance_0054 <= 920306;
    i_distance_0055 <= 845683;
    i_distance_0056 <= 48626;
    i_distance_0057 <= 404725;
    i_distance_0058 <= 142326;
    i_distance_0059 <= 303859;
    i_distance_0060 <= 485618;
    i_distance_0061 <= 1008757;
    i_distance_0062 <= 377466;
    i_distance_0063 <= 477947;
    correct_answer <= 15884;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 833921;
    i_distance_0001 <= 1005570;
    i_distance_0002 <= 785411;
    i_distance_0003 <= 394244;
    i_distance_0004 <= 177288;
    i_distance_0005 <= 414346;
    i_distance_0006 <= 587018;
    i_distance_0007 <= 175756;
    i_distance_0008 <= 764943;
    i_distance_0009 <= 430607;
    i_distance_0010 <= 948498;
    i_distance_0011 <= 267672;
    i_distance_0012 <= 594585;
    i_distance_0013 <= 60184;
    i_distance_0014 <= 537371;
    i_distance_0015 <= 835617;
    i_distance_0016 <= 255395;
    i_distance_0017 <= 964260;
    i_distance_0018 <= 98340;
    i_distance_0019 <= 171046;
    i_distance_0020 <= 166312;
    i_distance_0021 <= 366636;
    i_distance_0022 <= 917423;
    i_distance_0023 <= 530866;
    i_distance_0024 <= 767027;
    i_distance_0025 <= 630836;
    i_distance_0026 <= 148532;
    i_distance_0027 <= 234679;
    i_distance_0028 <= 365751;
    i_distance_0029 <= 903351;
    i_distance_0030 <= 436223;
    i_distance_0031 <= 264124;
    i_distance_0032 <= 901565;
    i_distance_0033 <= 819134;
    i_distance_0034 <= 65598;
    i_distance_0035 <= 578752;
    i_distance_0036 <= 869820;
    i_distance_0037 <= 373314;
    i_distance_0038 <= 679618;
    i_distance_0039 <= 640452;
    i_distance_0040 <= 449604;
    i_distance_0041 <= 624070;
    i_distance_0042 <= 601415;
    i_distance_0043 <= 96841;
    i_distance_0044 <= 760138;
    i_distance_0045 <= 340553;
    i_distance_0046 <= 5836;
    i_distance_0047 <= 111949;
    i_distance_0048 <= 805709;
    i_distance_0049 <= 886349;
    i_distance_0050 <= 526287;
    i_distance_0051 <= 97619;
    i_distance_0052 <= 648916;
    i_distance_0053 <= 431198;
    i_distance_0054 <= 646757;
    i_distance_0055 <= 313189;
    i_distance_0056 <= 560619;
    i_distance_0057 <= 924779;
    i_distance_0058 <= 1009775;
    i_distance_0059 <= 440176;
    i_distance_0060 <= 659188;
    i_distance_0061 <= 82932;
    i_distance_0062 <= 559227;
    i_distance_0063 <= 135679;
    correct_answer <= 5836;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 172161;
    i_distance_0001 <= 386561;
    i_distance_0002 <= 227334;
    i_distance_0003 <= 55815;
    i_distance_0004 <= 626056;
    i_distance_0005 <= 414857;
    i_distance_0006 <= 390923;
    i_distance_0007 <= 508174;
    i_distance_0008 <= 303122;
    i_distance_0009 <= 63763;
    i_distance_0010 <= 239765;
    i_distance_0011 <= 192409;
    i_distance_0012 <= 108953;
    i_distance_0013 <= 15385;
    i_distance_0014 <= 431006;
    i_distance_0015 <= 473759;
    i_distance_0016 <= 366497;
    i_distance_0017 <= 684069;
    i_distance_0018 <= 433959;
    i_distance_0019 <= 344233;
    i_distance_0020 <= 649514;
    i_distance_0021 <= 228394;
    i_distance_0022 <= 219180;
    i_distance_0023 <= 388522;
    i_distance_0024 <= 658736;
    i_distance_0025 <= 355120;
    i_distance_0026 <= 517682;
    i_distance_0027 <= 542258;
    i_distance_0028 <= 400690;
    i_distance_0029 <= 893371;
    i_distance_0030 <= 656956;
    i_distance_0031 <= 485819;
    i_distance_0032 <= 641853;
    i_distance_0033 <= 903999;
    i_distance_0034 <= 140608;
    i_distance_0035 <= 682308;
    i_distance_0036 <= 153032;
    i_distance_0037 <= 714441;
    i_distance_0038 <= 135246;
    i_distance_0039 <= 199887;
    i_distance_0040 <= 93134;
    i_distance_0041 <= 795985;
    i_distance_0042 <= 733135;
    i_distance_0043 <= 699605;
    i_distance_0044 <= 48214;
    i_distance_0045 <= 875861;
    i_distance_0046 <= 760026;
    i_distance_0047 <= 897374;
    i_distance_0048 <= 709471;
    i_distance_0049 <= 607848;
    i_distance_0050 <= 824425;
    i_distance_0051 <= 920298;
    i_distance_0052 <= 703720;
    i_distance_0053 <= 882670;
    i_distance_0054 <= 456303;
    i_distance_0055 <= 723566;
    i_distance_0056 <= 46703;
    i_distance_0057 <= 815854;
    i_distance_0058 <= 630131;
    i_distance_0059 <= 89460;
    i_distance_0060 <= 770166;
    i_distance_0061 <= 837110;
    i_distance_0062 <= 491256;
    i_distance_0063 <= 992123;
    correct_answer <= 15385;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 431362;
    i_distance_0001 <= 849411;
    i_distance_0002 <= 762498;
    i_distance_0003 <= 857735;
    i_distance_0004 <= 73480;
    i_distance_0005 <= 357387;
    i_distance_0006 <= 357004;
    i_distance_0007 <= 1032081;
    i_distance_0008 <= 110995;
    i_distance_0009 <= 434324;
    i_distance_0010 <= 685945;
    i_distance_0011 <= 503834;
    i_distance_0012 <= 776092;
    i_distance_0013 <= 979616;
    i_distance_0014 <= 725666;
    i_distance_0015 <= 421414;
    i_distance_0016 <= 602410;
    i_distance_0017 <= 504234;
    i_distance_0018 <= 627758;
    i_distance_0019 <= 485553;
    i_distance_0020 <= 631858;
    i_distance_0021 <= 1033397;
    i_distance_0022 <= 798775;
    i_distance_0023 <= 20537;
    i_distance_0024 <= 79806;
    i_distance_0025 <= 525758;
    i_distance_0026 <= 268863;
    i_distance_0027 <= 955198;
    i_distance_0028 <= 991171;
    i_distance_0029 <= 424390;
    i_distance_0030 <= 346696;
    i_distance_0031 <= 147785;
    i_distance_0032 <= 362314;
    i_distance_0033 <= 237258;
    i_distance_0034 <= 634190;
    i_distance_0035 <= 498513;
    i_distance_0036 <= 667258;
    i_distance_0037 <= 10072;
    i_distance_0038 <= 438363;
    i_distance_0039 <= 365918;
    i_distance_0040 <= 264032;
    i_distance_0041 <= 104929;
    i_distance_0042 <= 456160;
    i_distance_0043 <= 608355;
    i_distance_0044 <= 979297;
    i_distance_0045 <= 42608;
    i_distance_0046 <= 295016;
    i_distance_0047 <= 953580;
    i_distance_0048 <= 492781;
    i_distance_0049 <= 380911;
    i_distance_0050 <= 593392;
    i_distance_0051 <= 28913;
    i_distance_0052 <= 117618;
    i_distance_0053 <= 74355;
    i_distance_0054 <= 96884;
    i_distance_0055 <= 774640;
    i_distance_0056 <= 141686;
    i_distance_0057 <= 966903;
    i_distance_0058 <= 439160;
    i_distance_0059 <= 836344;
    i_distance_0060 <= 452213;
    i_distance_0061 <= 440955;
    i_distance_0062 <= 3196;
    i_distance_0063 <= 986367;
    correct_answer <= 3196;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 449798;
    i_distance_0001 <= 531206;
    i_distance_0002 <= 503305;
    i_distance_0003 <= 682762;
    i_distance_0004 <= 296971;
    i_distance_0005 <= 972298;
    i_distance_0006 <= 199564;
    i_distance_0007 <= 731019;
    i_distance_0008 <= 344585;
    i_distance_0009 <= 279060;
    i_distance_0010 <= 649493;
    i_distance_0011 <= 267669;
    i_distance_0012 <= 954136;
    i_distance_0013 <= 145433;
    i_distance_0014 <= 885403;
    i_distance_0015 <= 444187;
    i_distance_0016 <= 66077;
    i_distance_0017 <= 718878;
    i_distance_0018 <= 318369;
    i_distance_0019 <= 674594;
    i_distance_0020 <= 492195;
    i_distance_0021 <= 255907;
    i_distance_0022 <= 766375;
    i_distance_0023 <= 1040040;
    i_distance_0024 <= 947115;
    i_distance_0025 <= 563372;
    i_distance_0026 <= 642992;
    i_distance_0027 <= 744374;
    i_distance_0028 <= 1042233;
    i_distance_0029 <= 379840;
    i_distance_0030 <= 695745;
    i_distance_0031 <= 1007552;
    i_distance_0032 <= 79171;
    i_distance_0033 <= 531396;
    i_distance_0034 <= 280267;
    i_distance_0035 <= 354379;
    i_distance_0036 <= 344017;
    i_distance_0037 <= 987474;
    i_distance_0038 <= 727505;
    i_distance_0039 <= 286932;
    i_distance_0040 <= 136917;
    i_distance_0041 <= 1001688;
    i_distance_0042 <= 363357;
    i_distance_0043 <= 651615;
    i_distance_0044 <= 489697;
    i_distance_0045 <= 443363;
    i_distance_0046 <= 210277;
    i_distance_0047 <= 274664;
    i_distance_0048 <= 452329;
    i_distance_0049 <= 173289;
    i_distance_0050 <= 24171;
    i_distance_0051 <= 965611;
    i_distance_0052 <= 343788;
    i_distance_0053 <= 842736;
    i_distance_0054 <= 450928;
    i_distance_0055 <= 62835;
    i_distance_0056 <= 950900;
    i_distance_0057 <= 354549;
    i_distance_0058 <= 353142;
    i_distance_0059 <= 549496;
    i_distance_0060 <= 157305;
    i_distance_0061 <= 97531;
    i_distance_0062 <= 390142;
    i_distance_0063 <= 74495;
    correct_answer <= 24171;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 853760;
    i_distance_0001 <= 103425;
    i_distance_0002 <= 140417;
    i_distance_0003 <= 744705;
    i_distance_0004 <= 676226;
    i_distance_0005 <= 181637;
    i_distance_0006 <= 357896;
    i_distance_0007 <= 243208;
    i_distance_0008 <= 316298;
    i_distance_0009 <= 392842;
    i_distance_0010 <= 145932;
    i_distance_0011 <= 101005;
    i_distance_0012 <= 678029;
    i_distance_0013 <= 501138;
    i_distance_0014 <= 82450;
    i_distance_0015 <= 994969;
    i_distance_0016 <= 477210;
    i_distance_0017 <= 243611;
    i_distance_0018 <= 257566;
    i_distance_0019 <= 463649;
    i_distance_0020 <= 522916;
    i_distance_0021 <= 900516;
    i_distance_0022 <= 2214;
    i_distance_0023 <= 114349;
    i_distance_0024 <= 173104;
    i_distance_0025 <= 190516;
    i_distance_0026 <= 396085;
    i_distance_0027 <= 5942;
    i_distance_0028 <= 740791;
    i_distance_0029 <= 728757;
    i_distance_0030 <= 10806;
    i_distance_0031 <= 705850;
    i_distance_0032 <= 613303;
    i_distance_0033 <= 350079;
    i_distance_0034 <= 159417;
    i_distance_0035 <= 389953;
    i_distance_0036 <= 838084;
    i_distance_0037 <= 335813;
    i_distance_0038 <= 1030086;
    i_distance_0039 <= 784840;
    i_distance_0040 <= 652877;
    i_distance_0041 <= 1003726;
    i_distance_0042 <= 882259;
    i_distance_0043 <= 102106;
    i_distance_0044 <= 933723;
    i_distance_0045 <= 173150;
    i_distance_0046 <= 176611;
    i_distance_0047 <= 381924;
    i_distance_0048 <= 851686;
    i_distance_0049 <= 950631;
    i_distance_0050 <= 423911;
    i_distance_0051 <= 776425;
    i_distance_0052 <= 704620;
    i_distance_0053 <= 1034861;
    i_distance_0054 <= 880494;
    i_distance_0055 <= 578797;
    i_distance_0056 <= 644973;
    i_distance_0057 <= 776428;
    i_distance_0058 <= 947186;
    i_distance_0059 <= 944243;
    i_distance_0060 <= 164472;
    i_distance_0061 <= 806393;
    i_distance_0062 <= 511486;
    i_distance_0063 <= 348415;
    correct_answer <= 2214;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 753920;
    i_distance_0001 <= 176386;
    i_distance_0002 <= 356354;
    i_distance_0003 <= 282630;
    i_distance_0004 <= 33158;
    i_distance_0005 <= 648073;
    i_distance_0006 <= 1032202;
    i_distance_0007 <= 300555;
    i_distance_0008 <= 641545;
    i_distance_0009 <= 761740;
    i_distance_0010 <= 930190;
    i_distance_0011 <= 33042;
    i_distance_0012 <= 14995;
    i_distance_0013 <= 616340;
    i_distance_0014 <= 458389;
    i_distance_0015 <= 688146;
    i_distance_0016 <= 410142;
    i_distance_0017 <= 492063;
    i_distance_0018 <= 26109;
    i_distance_0019 <= 707747;
    i_distance_0020 <= 967847;
    i_distance_0021 <= 971305;
    i_distance_0022 <= 306351;
    i_distance_0023 <= 718640;
    i_distance_0024 <= 162225;
    i_distance_0025 <= 269617;
    i_distance_0026 <= 216117;
    i_distance_0027 <= 726584;
    i_distance_0028 <= 800824;
    i_distance_0029 <= 198328;
    i_distance_0030 <= 511424;
    i_distance_0031 <= 404289;
    i_distance_0032 <= 543042;
    i_distance_0033 <= 305732;
    i_distance_0034 <= 596293;
    i_distance_0035 <= 777925;
    i_distance_0036 <= 22598;
    i_distance_0037 <= 74824;
    i_distance_0038 <= 848200;
    i_distance_0039 <= 50628;
    i_distance_0040 <= 302925;
    i_distance_0041 <= 653008;
    i_distance_0042 <= 1004242;
    i_distance_0043 <= 798675;
    i_distance_0044 <= 674260;
    i_distance_0045 <= 81748;
    i_distance_0046 <= 388181;
    i_distance_0047 <= 166875;
    i_distance_0048 <= 285917;
    i_distance_0049 <= 580833;
    i_distance_0050 <= 286050;
    i_distance_0051 <= 65251;
    i_distance_0052 <= 755435;
    i_distance_0053 <= 68974;
    i_distance_0054 <= 96111;
    i_distance_0055 <= 221939;
    i_distance_0056 <= 102779;
    i_distance_0057 <= 165622;
    i_distance_0058 <= 430583;
    i_distance_0059 <= 534008;
    i_distance_0060 <= 745850;
    i_distance_0061 <= 174587;
    i_distance_0062 <= 686716;
    i_distance_0063 <= 221949;
    correct_answer <= 14995;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 836984;
    i_distance_0001 <= 719620;
    i_distance_0002 <= 555784;
    i_distance_0003 <= 491528;
    i_distance_0004 <= 198411;
    i_distance_0005 <= 684939;
    i_distance_0006 <= 817420;
    i_distance_0007 <= 700435;
    i_distance_0008 <= 630932;
    i_distance_0009 <= 12691;
    i_distance_0010 <= 1046934;
    i_distance_0011 <= 312954;
    i_distance_0012 <= 256156;
    i_distance_0013 <= 651293;
    i_distance_0014 <= 192030;
    i_distance_0015 <= 482721;
    i_distance_0016 <= 285091;
    i_distance_0017 <= 425635;
    i_distance_0018 <= 720421;
    i_distance_0019 <= 635050;
    i_distance_0020 <= 721964;
    i_distance_0021 <= 833328;
    i_distance_0022 <= 312881;
    i_distance_0023 <= 945202;
    i_distance_0024 <= 108857;
    i_distance_0025 <= 634428;
    i_distance_0026 <= 714557;
    i_distance_0027 <= 947910;
    i_distance_0028 <= 355661;
    i_distance_0029 <= 20302;
    i_distance_0030 <= 662736;
    i_distance_0031 <= 483281;
    i_distance_0032 <= 814034;
    i_distance_0033 <= 836819;
    i_distance_0034 <= 179030;
    i_distance_0035 <= 111703;
    i_distance_0036 <= 809432;
    i_distance_0037 <= 493656;
    i_distance_0038 <= 64728;
    i_distance_0039 <= 261849;
    i_distance_0040 <= 534239;
    i_distance_0041 <= 447712;
    i_distance_0042 <= 374498;
    i_distance_0043 <= 16100;
    i_distance_0044 <= 454503;
    i_distance_0045 <= 367336;
    i_distance_0046 <= 638057;
    i_distance_0047 <= 748905;
    i_distance_0048 <= 87275;
    i_distance_0049 <= 403052;
    i_distance_0050 <= 803308;
    i_distance_0051 <= 593646;
    i_distance_0052 <= 837487;
    i_distance_0053 <= 399856;
    i_distance_0054 <= 904049;
    i_distance_0055 <= 442874;
    i_distance_0056 <= 193514;
    i_distance_0057 <= 374134;
    i_distance_0058 <= 226678;
    i_distance_0059 <= 671096;
    i_distance_0060 <= 903034;
    i_distance_0061 <= 1040507;
    i_distance_0062 <= 294397;
    i_distance_0063 <= 189311;
    correct_answer <= 12691;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 402949;
    i_distance_0001 <= 101640;
    i_distance_0002 <= 509448;
    i_distance_0003 <= 964108;
    i_distance_0004 <= 294797;
    i_distance_0005 <= 561038;
    i_distance_0006 <= 264081;
    i_distance_0007 <= 112785;
    i_distance_0008 <= 371860;
    i_distance_0009 <= 11541;
    i_distance_0010 <= 780951;
    i_distance_0011 <= 112408;
    i_distance_0012 <= 330650;
    i_distance_0013 <= 88218;
    i_distance_0014 <= 904220;
    i_distance_0015 <= 499490;
    i_distance_0016 <= 686882;
    i_distance_0017 <= 591397;
    i_distance_0018 <= 665128;
    i_distance_0019 <= 712106;
    i_distance_0020 <= 1048107;
    i_distance_0021 <= 5804;
    i_distance_0022 <= 252973;
    i_distance_0023 <= 643374;
    i_distance_0024 <= 55470;
    i_distance_0025 <= 622766;
    i_distance_0026 <= 260657;
    i_distance_0027 <= 505651;
    i_distance_0028 <= 326837;
    i_distance_0029 <= 673078;
    i_distance_0030 <= 854843;
    i_distance_0031 <= 829117;
    i_distance_0032 <= 436159;
    i_distance_0033 <= 402239;
    i_distance_0034 <= 778945;
    i_distance_0035 <= 189507;
    i_distance_0036 <= 953028;
    i_distance_0037 <= 197575;
    i_distance_0038 <= 266314;
    i_distance_0039 <= 58442;
    i_distance_0040 <= 312396;
    i_distance_0041 <= 536397;
    i_distance_0042 <= 839630;
    i_distance_0043 <= 654548;
    i_distance_0044 <= 804052;
    i_distance_0045 <= 885076;
    i_distance_0046 <= 265431;
    i_distance_0047 <= 563416;
    i_distance_0048 <= 42967;
    i_distance_0049 <= 292181;
    i_distance_0050 <= 760545;
    i_distance_0051 <= 489955;
    i_distance_0052 <= 719716;
    i_distance_0053 <= 348131;
    i_distance_0054 <= 767204;
    i_distance_0055 <= 852198;
    i_distance_0056 <= 48746;
    i_distance_0057 <= 536690;
    i_distance_0058 <= 509555;
    i_distance_0059 <= 89076;
    i_distance_0060 <= 308855;
    i_distance_0061 <= 903800;
    i_distance_0062 <= 470521;
    i_distance_0063 <= 696314;
    correct_answer <= 5804;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 890627;
    i_distance_0001 <= 857348;
    i_distance_0002 <= 524166;
    i_distance_0003 <= 126856;
    i_distance_0004 <= 233998;
    i_distance_0005 <= 534286;
    i_distance_0006 <= 441493;
    i_distance_0007 <= 1039254;
    i_distance_0008 <= 397975;
    i_distance_0009 <= 589079;
    i_distance_0010 <= 280984;
    i_distance_0011 <= 359450;
    i_distance_0012 <= 870170;
    i_distance_0013 <= 91676;
    i_distance_0014 <= 123933;
    i_distance_0015 <= 1019038;
    i_distance_0016 <= 653858;
    i_distance_0017 <= 889764;
    i_distance_0018 <= 1039653;
    i_distance_0019 <= 771366;
    i_distance_0020 <= 930987;
    i_distance_0021 <= 479149;
    i_distance_0022 <= 783917;
    i_distance_0023 <= 905647;
    i_distance_0024 <= 268847;
    i_distance_0025 <= 577074;
    i_distance_0026 <= 140597;
    i_distance_0027 <= 68662;
    i_distance_0028 <= 107703;
    i_distance_0029 <= 871099;
    i_distance_0030 <= 1002428;
    i_distance_0031 <= 908860;
    i_distance_0032 <= 1019201;
    i_distance_0033 <= 290370;
    i_distance_0034 <= 971585;
    i_distance_0035 <= 552513;
    i_distance_0036 <= 665925;
    i_distance_0037 <= 155461;
    i_distance_0038 <= 883525;
    i_distance_0039 <= 222794;
    i_distance_0040 <= 117578;
    i_distance_0041 <= 436815;
    i_distance_0042 <= 197073;
    i_distance_0043 <= 964181;
    i_distance_0044 <= 769242;
    i_distance_0045 <= 317532;
    i_distance_0046 <= 44509;
    i_distance_0047 <= 756061;
    i_distance_0048 <= 471133;
    i_distance_0049 <= 544352;
    i_distance_0050 <= 893154;
    i_distance_0051 <= 32867;
    i_distance_0052 <= 100067;
    i_distance_0053 <= 890724;
    i_distance_0054 <= 662883;
    i_distance_0055 <= 241895;
    i_distance_0056 <= 1026922;
    i_distance_0057 <= 464618;
    i_distance_0058 <= 830058;
    i_distance_0059 <= 392436;
    i_distance_0060 <= 427637;
    i_distance_0061 <= 168184;
    i_distance_0062 <= 556028;
    i_distance_0063 <= 693245;
    correct_answer <= 32867;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 117763;
    i_distance_0001 <= 94084;
    i_distance_0002 <= 743432;
    i_distance_0003 <= 394890;
    i_distance_0004 <= 193419;
    i_distance_0005 <= 780300;
    i_distance_0006 <= 840719;
    i_distance_0007 <= 1032594;
    i_distance_0008 <= 118802;
    i_distance_0009 <= 185748;
    i_distance_0010 <= 27412;
    i_distance_0011 <= 290965;
    i_distance_0012 <= 1037591;
    i_distance_0013 <= 535576;
    i_distance_0014 <= 171549;
    i_distance_0015 <= 1042339;
    i_distance_0016 <= 274851;
    i_distance_0017 <= 6693;
    i_distance_0018 <= 751908;
    i_distance_0019 <= 634916;
    i_distance_0020 <= 58281;
    i_distance_0021 <= 698538;
    i_distance_0022 <= 969131;
    i_distance_0023 <= 836525;
    i_distance_0024 <= 901424;
    i_distance_0025 <= 824625;
    i_distance_0026 <= 210226;
    i_distance_0027 <= 1025331;
    i_distance_0028 <= 305460;
    i_distance_0029 <= 609971;
    i_distance_0030 <= 965556;
    i_distance_0031 <= 379700;
    i_distance_0032 <= 213944;
    i_distance_0033 <= 89657;
    i_distance_0034 <= 709946;
    i_distance_0035 <= 854209;
    i_distance_0036 <= 972226;
    i_distance_0037 <= 331202;
    i_distance_0038 <= 535491;
    i_distance_0039 <= 1036355;
    i_distance_0040 <= 418499;
    i_distance_0041 <= 856898;
    i_distance_0042 <= 578376;
    i_distance_0043 <= 272713;
    i_distance_0044 <= 325062;
    i_distance_0045 <= 622923;
    i_distance_0046 <= 529996;
    i_distance_0047 <= 759626;
    i_distance_0048 <= 449612;
    i_distance_0049 <= 398800;
    i_distance_0050 <= 619358;
    i_distance_0051 <= 216828;
    i_distance_0052 <= 298984;
    i_distance_0053 <= 57832;
    i_distance_0054 <= 393960;
    i_distance_0055 <= 916207;
    i_distance_0056 <= 432625;
    i_distance_0057 <= 166386;
    i_distance_0058 <= 511221;
    i_distance_0059 <= 618358;
    i_distance_0060 <= 510455;
    i_distance_0061 <= 841850;
    i_distance_0062 <= 721147;
    i_distance_0063 <= 96636;
    correct_answer <= 6693;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 100865;
    i_distance_0001 <= 772231;
    i_distance_0002 <= 349064;
    i_distance_0003 <= 354184;
    i_distance_0004 <= 335117;
    i_distance_0005 <= 70542;
    i_distance_0006 <= 320400;
    i_distance_0007 <= 895637;
    i_distance_0008 <= 570008;
    i_distance_0009 <= 447258;
    i_distance_0010 <= 905756;
    i_distance_0011 <= 992285;
    i_distance_0012 <= 489246;
    i_distance_0013 <= 928542;
    i_distance_0014 <= 882976;
    i_distance_0015 <= 481821;
    i_distance_0016 <= 514424;
    i_distance_0017 <= 726437;
    i_distance_0018 <= 210344;
    i_distance_0019 <= 862248;
    i_distance_0020 <= 1030959;
    i_distance_0021 <= 514097;
    i_distance_0022 <= 906804;
    i_distance_0023 <= 384059;
    i_distance_0024 <= 880317;
    i_distance_0025 <= 781501;
    i_distance_0026 <= 4161;
    i_distance_0027 <= 860099;
    i_distance_0028 <= 929735;
    i_distance_0029 <= 103496;
    i_distance_0030 <= 904266;
    i_distance_0031 <= 302539;
    i_distance_0032 <= 452172;
    i_distance_0033 <= 849740;
    i_distance_0034 <= 116554;
    i_distance_0035 <= 138321;
    i_distance_0036 <= 454356;
    i_distance_0037 <= 558679;
    i_distance_0038 <= 631000;
    i_distance_0039 <= 873945;
    i_distance_0040 <= 742493;
    i_distance_0041 <= 663392;
    i_distance_0042 <= 562529;
    i_distance_0043 <= 61410;
    i_distance_0044 <= 551523;
    i_distance_0045 <= 229604;
    i_distance_0046 <= 111589;
    i_distance_0047 <= 383206;
    i_distance_0048 <= 21478;
    i_distance_0049 <= 1022692;
    i_distance_0050 <= 186089;
    i_distance_0051 <= 842090;
    i_distance_0052 <= 671852;
    i_distance_0053 <= 44270;
    i_distance_0054 <= 937328;
    i_distance_0055 <= 392048;
    i_distance_0056 <= 99443;
    i_distance_0057 <= 775669;
    i_distance_0058 <= 899829;
    i_distance_0059 <= 397429;
    i_distance_0060 <= 287224;
    i_distance_0061 <= 900730;
    i_distance_0062 <= 884219;
    i_distance_0063 <= 710653;
    correct_answer <= 4161;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 352386;
    i_distance_0001 <= 888452;
    i_distance_0002 <= 79493;
    i_distance_0003 <= 670856;
    i_distance_0004 <= 540041;
    i_distance_0005 <= 912524;
    i_distance_0006 <= 1040270;
    i_distance_0007 <= 1042576;
    i_distance_0008 <= 134162;
    i_distance_0009 <= 947986;
    i_distance_0010 <= 360467;
    i_distance_0011 <= 404886;
    i_distance_0012 <= 268695;
    i_distance_0013 <= 162586;
    i_distance_0014 <= 386333;
    i_distance_0015 <= 500770;
    i_distance_0016 <= 47907;
    i_distance_0017 <= 963966;
    i_distance_0018 <= 31911;
    i_distance_0019 <= 287530;
    i_distance_0020 <= 280236;
    i_distance_0021 <= 420911;
    i_distance_0022 <= 783279;
    i_distance_0023 <= 744496;
    i_distance_0024 <= 444340;
    i_distance_0025 <= 606260;
    i_distance_0026 <= 114613;
    i_distance_0027 <= 770361;
    i_distance_0028 <= 419258;
    i_distance_0029 <= 649659;
    i_distance_0030 <= 615100;
    i_distance_0031 <= 115901;
    i_distance_0032 <= 629821;
    i_distance_0033 <= 320062;
    i_distance_0034 <= 887739;
    i_distance_0035 <= 604091;
    i_distance_0036 <= 504768;
    i_distance_0037 <= 966725;
    i_distance_0038 <= 795207;
    i_distance_0039 <= 564808;
    i_distance_0040 <= 93383;
    i_distance_0041 <= 914254;
    i_distance_0042 <= 657617;
    i_distance_0043 <= 881746;
    i_distance_0044 <= 155091;
    i_distance_0045 <= 974676;
    i_distance_0046 <= 591958;
    i_distance_0047 <= 776409;
    i_distance_0048 <= 441182;
    i_distance_0049 <= 31584;
    i_distance_0050 <= 771680;
    i_distance_0051 <= 135909;
    i_distance_0052 <= 1045863;
    i_distance_0053 <= 71271;
    i_distance_0054 <= 689386;
    i_distance_0055 <= 451821;
    i_distance_0056 <= 643821;
    i_distance_0057 <= 645231;
    i_distance_0058 <= 422000;
    i_distance_0059 <= 420596;
    i_distance_0060 <= 388469;
    i_distance_0061 <= 303349;
    i_distance_0062 <= 861559;
    i_distance_0063 <= 94206;
    correct_answer <= 31584;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 82304;
    i_distance_0001 <= 37380;
    i_distance_0002 <= 34693;
    i_distance_0003 <= 590340;
    i_distance_0004 <= 602245;
    i_distance_0005 <= 518409;
    i_distance_0006 <= 242825;
    i_distance_0007 <= 31370;
    i_distance_0008 <= 620429;
    i_distance_0009 <= 769553;
    i_distance_0010 <= 665618;
    i_distance_0011 <= 155544;
    i_distance_0012 <= 207514;
    i_distance_0013 <= 696090;
    i_distance_0014 <= 286620;
    i_distance_0015 <= 654877;
    i_distance_0016 <= 328480;
    i_distance_0017 <= 493857;
    i_distance_0018 <= 951466;
    i_distance_0019 <= 805932;
    i_distance_0020 <= 682924;
    i_distance_0021 <= 523951;
    i_distance_0022 <= 702768;
    i_distance_0023 <= 138801;
    i_distance_0024 <= 999475;
    i_distance_0025 <= 875827;
    i_distance_0026 <= 284213;
    i_distance_0027 <= 441397;
    i_distance_0028 <= 1041717;
    i_distance_0029 <= 599608;
    i_distance_0030 <= 921782;
    i_distance_0031 <= 914752;
    i_distance_0032 <= 709953;
    i_distance_0033 <= 326464;
    i_distance_0034 <= 34115;
    i_distance_0035 <= 423364;
    i_distance_0036 <= 574784;
    i_distance_0037 <= 449991;
    i_distance_0038 <= 977224;
    i_distance_0039 <= 1035211;
    i_distance_0040 <= 820945;
    i_distance_0041 <= 704978;
    i_distance_0042 <= 871125;
    i_distance_0043 <= 911958;
    i_distance_0044 <= 690007;
    i_distance_0045 <= 765401;
    i_distance_0046 <= 382297;
    i_distance_0047 <= 1020124;
    i_distance_0048 <= 716128;
    i_distance_0049 <= 594662;
    i_distance_0050 <= 342503;
    i_distance_0051 <= 988521;
    i_distance_0052 <= 545641;
    i_distance_0053 <= 537962;
    i_distance_0054 <= 659565;
    i_distance_0055 <= 922990;
    i_distance_0056 <= 383727;
    i_distance_0057 <= 431477;
    i_distance_0058 <= 977910;
    i_distance_0059 <= 187383;
    i_distance_0060 <= 106617;
    i_distance_0061 <= 587002;
    i_distance_0062 <= 986109;
    i_distance_0063 <= 233599;
    correct_answer <= 31370;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 615040;
    i_distance_0001 <= 12033;
    i_distance_0002 <= 179074;
    i_distance_0003 <= 165252;
    i_distance_0004 <= 860677;
    i_distance_0005 <= 142728;
    i_distance_0006 <= 424201;
    i_distance_0007 <= 451467;
    i_distance_0008 <= 401036;
    i_distance_0009 <= 148222;
    i_distance_0010 <= 739600;
    i_distance_0011 <= 741904;
    i_distance_0012 <= 419090;
    i_distance_0013 <= 60432;
    i_distance_0014 <= 313876;
    i_distance_0015 <= 7701;
    i_distance_0016 <= 361752;
    i_distance_0017 <= 53656;
    i_distance_0018 <= 940826;
    i_distance_0019 <= 1034524;
    i_distance_0020 <= 459037;
    i_distance_0021 <= 653216;
    i_distance_0022 <= 993443;
    i_distance_0023 <= 814118;
    i_distance_0024 <= 494886;
    i_distance_0025 <= 505896;
    i_distance_0026 <= 192038;
    i_distance_0027 <= 838954;
    i_distance_0028 <= 600620;
    i_distance_0029 <= 324908;
    i_distance_0030 <= 983214;
    i_distance_0031 <= 186170;
    i_distance_0032 <= 1033408;
    i_distance_0033 <= 141761;
    i_distance_0034 <= 876864;
    i_distance_0035 <= 972486;
    i_distance_0036 <= 874439;
    i_distance_0037 <= 745287;
    i_distance_0038 <= 162763;
    i_distance_0039 <= 151628;
    i_distance_0040 <= 406861;
    i_distance_0041 <= 138573;
    i_distance_0042 <= 365774;
    i_distance_0043 <= 806478;
    i_distance_0044 <= 322895;
    i_distance_0045 <= 804561;
    i_distance_0046 <= 229719;
    i_distance_0047 <= 264407;
    i_distance_0048 <= 968153;
    i_distance_0049 <= 30810;
    i_distance_0050 <= 1014103;
    i_distance_0051 <= 664924;
    i_distance_0052 <= 79583;
    i_distance_0053 <= 715233;
    i_distance_0054 <= 315237;
    i_distance_0055 <= 843367;
    i_distance_0056 <= 326249;
    i_distance_0057 <= 143465;
    i_distance_0058 <= 758895;
    i_distance_0059 <= 153072;
    i_distance_0060 <= 1006706;
    i_distance_0061 <= 863990;
    i_distance_0062 <= 744958;
    i_distance_0063 <= 912639;
    correct_answer <= 7701;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 218498;
    i_distance_0001 <= 1029380;
    i_distance_0002 <= 308870;
    i_distance_0003 <= 809095;
    i_distance_0004 <= 915335;
    i_distance_0005 <= 272394;
    i_distance_0006 <= 537723;
    i_distance_0007 <= 869520;
    i_distance_0008 <= 35216;
    i_distance_0009 <= 1035027;
    i_distance_0010 <= 120086;
    i_distance_0011 <= 867738;
    i_distance_0012 <= 928411;
    i_distance_0013 <= 242076;
    i_distance_0014 <= 835226;
    i_distance_0015 <= 339485;
    i_distance_0016 <= 419871;
    i_distance_0017 <= 968609;
    i_distance_0018 <= 200738;
    i_distance_0019 <= 317606;
    i_distance_0020 <= 607783;
    i_distance_0021 <= 444073;
    i_distance_0022 <= 17450;
    i_distance_0023 <= 74156;
    i_distance_0024 <= 125306;
    i_distance_0025 <= 292399;
    i_distance_0026 <= 330545;
    i_distance_0027 <= 347827;
    i_distance_0028 <= 363130;
    i_distance_0029 <= 271801;
    i_distance_0030 <= 313146;
    i_distance_0031 <= 367036;
    i_distance_0032 <= 581058;
    i_distance_0033 <= 17476;
    i_distance_0034 <= 123460;
    i_distance_0035 <= 1038793;
    i_distance_0036 <= 509514;
    i_distance_0037 <= 461387;
    i_distance_0038 <= 823625;
    i_distance_0039 <= 576846;
    i_distance_0040 <= 626895;
    i_distance_0041 <= 124625;
    i_distance_0042 <= 747347;
    i_distance_0043 <= 409719;
    i_distance_0044 <= 984539;
    i_distance_0045 <= 978810;
    i_distance_0046 <= 568415;
    i_distance_0047 <= 243552;
    i_distance_0048 <= 715232;
    i_distance_0049 <= 918883;
    i_distance_0050 <= 189158;
    i_distance_0051 <= 270568;
    i_distance_0052 <= 824554;
    i_distance_0053 <= 834795;
    i_distance_0054 <= 671725;
    i_distance_0055 <= 894447;
    i_distance_0056 <= 39279;
    i_distance_0057 <= 291953;
    i_distance_0058 <= 979826;
    i_distance_0059 <= 379767;
    i_distance_0060 <= 25850;
    i_distance_0061 <= 9339;
    i_distance_0062 <= 4476;
    i_distance_0063 <= 434175;
    correct_answer <= 4476;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 666629;
    i_distance_0001 <= 338566;
    i_distance_0002 <= 1003658;
    i_distance_0003 <= 361867;
    i_distance_0004 <= 585490;
    i_distance_0005 <= 243347;
    i_distance_0006 <= 215828;
    i_distance_0007 <= 521112;
    i_distance_0008 <= 1011612;
    i_distance_0009 <= 225184;
    i_distance_0010 <= 587040;
    i_distance_0011 <= 669857;
    i_distance_0012 <= 731043;
    i_distance_0013 <= 836772;
    i_distance_0014 <= 453285;
    i_distance_0015 <= 973606;
    i_distance_0016 <= 12199;
    i_distance_0017 <= 857384;
    i_distance_0018 <= 133289;
    i_distance_0019 <= 617770;
    i_distance_0020 <= 846123;
    i_distance_0021 <= 575532;
    i_distance_0022 <= 251181;
    i_distance_0023 <= 978094;
    i_distance_0024 <= 662319;
    i_distance_0025 <= 170800;
    i_distance_0026 <= 303537;
    i_distance_0027 <= 491185;
    i_distance_0028 <= 136106;
    i_distance_0029 <= 914486;
    i_distance_0030 <= 221753;
    i_distance_0031 <= 820795;
    i_distance_0032 <= 4413;
    i_distance_0033 <= 834879;
    i_distance_0034 <= 716353;
    i_distance_0035 <= 410179;
    i_distance_0036 <= 681027;
    i_distance_0037 <= 845511;
    i_distance_0038 <= 893897;
    i_distance_0039 <= 951754;
    i_distance_0040 <= 473684;
    i_distance_0041 <= 369366;
    i_distance_0042 <= 1020023;
    i_distance_0043 <= 508632;
    i_distance_0044 <= 271704;
    i_distance_0045 <= 48598;
    i_distance_0046 <= 476383;
    i_distance_0047 <= 99554;
    i_distance_0048 <= 460130;
    i_distance_0049 <= 915684;
    i_distance_0050 <= 591083;
    i_distance_0051 <= 215020;
    i_distance_0052 <= 210797;
    i_distance_0053 <= 274285;
    i_distance_0054 <= 386287;
    i_distance_0055 <= 184689;
    i_distance_0056 <= 48754;
    i_distance_0057 <= 371956;
    i_distance_0058 <= 689398;
    i_distance_0059 <= 492791;
    i_distance_0060 <= 297848;
    i_distance_0061 <= 791930;
    i_distance_0062 <= 637949;
    i_distance_0063 <= 306686;
    correct_answer <= 4413;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 31361;
    i_distance_0001 <= 669579;
    i_distance_0002 <= 391054;
    i_distance_0003 <= 880655;
    i_distance_0004 <= 376850;
    i_distance_0005 <= 552467;
    i_distance_0006 <= 1026839;
    i_distance_0007 <= 532631;
    i_distance_0008 <= 256793;
    i_distance_0009 <= 889114;
    i_distance_0010 <= 455965;
    i_distance_0011 <= 148128;
    i_distance_0012 <= 453793;
    i_distance_0013 <= 480036;
    i_distance_0014 <= 247204;
    i_distance_0015 <= 530216;
    i_distance_0016 <= 970281;
    i_distance_0017 <= 340396;
    i_distance_0018 <= 360623;
    i_distance_0019 <= 105264;
    i_distance_0020 <= 516785;
    i_distance_0021 <= 876082;
    i_distance_0022 <= 984113;
    i_distance_0023 <= 436146;
    i_distance_0024 <= 819253;
    i_distance_0025 <= 629297;
    i_distance_0026 <= 42291;
    i_distance_0027 <= 331701;
    i_distance_0028 <= 211126;
    i_distance_0029 <= 271290;
    i_distance_0030 <= 595260;
    i_distance_0031 <= 823869;
    i_distance_0032 <= 576444;
    i_distance_0033 <= 828352;
    i_distance_0034 <= 989508;
    i_distance_0035 <= 915781;
    i_distance_0036 <= 299205;
    i_distance_0037 <= 89417;
    i_distance_0038 <= 773198;
    i_distance_0039 <= 485966;
    i_distance_0040 <= 819023;
    i_distance_0041 <= 108113;
    i_distance_0042 <= 810322;
    i_distance_0043 <= 115542;
    i_distance_0044 <= 688599;
    i_distance_0045 <= 738265;
    i_distance_0046 <= 393563;
    i_distance_0047 <= 72670;
    i_distance_0048 <= 701409;
    i_distance_0049 <= 957411;
    i_distance_0050 <= 25957;
    i_distance_0051 <= 320871;
    i_distance_0052 <= 429033;
    i_distance_0053 <= 137962;
    i_distance_0054 <= 1007211;
    i_distance_0055 <= 960620;
    i_distance_0056 <= 665325;
    i_distance_0057 <= 147568;
    i_distance_0058 <= 694005;
    i_distance_0059 <= 363383;
    i_distance_0060 <= 622456;
    i_distance_0061 <= 5625;
    i_distance_0062 <= 563194;
    i_distance_0063 <= 171644;
    correct_answer <= 5625;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 142723;
    i_distance_0001 <= 535556;
    i_distance_0002 <= 459014;
    i_distance_0003 <= 168583;
    i_distance_0004 <= 1027848;
    i_distance_0005 <= 996872;
    i_distance_0006 <= 57738;
    i_distance_0007 <= 868874;
    i_distance_0008 <= 109576;
    i_distance_0009 <= 65037;
    i_distance_0010 <= 963598;
    i_distance_0011 <= 1014163;
    i_distance_0012 <= 381973;
    i_distance_0013 <= 559893;
    i_distance_0014 <= 738199;
    i_distance_0015 <= 1020826;
    i_distance_0016 <= 514334;
    i_distance_0017 <= 246687;
    i_distance_0018 <= 728096;
    i_distance_0019 <= 714784;
    i_distance_0020 <= 167074;
    i_distance_0021 <= 182691;
    i_distance_0022 <= 934439;
    i_distance_0023 <= 377640;
    i_distance_0024 <= 82858;
    i_distance_0025 <= 327466;
    i_distance_0026 <= 580655;
    i_distance_0027 <= 530866;
    i_distance_0028 <= 406454;
    i_distance_0029 <= 786361;
    i_distance_0030 <= 525629;
    i_distance_0031 <= 846909;
    i_distance_0032 <= 582462;
    i_distance_0033 <= 633410;
    i_distance_0034 <= 986563;
    i_distance_0035 <= 807877;
    i_distance_0036 <= 720838;
    i_distance_0037 <= 651207;
    i_distance_0038 <= 809928;
    i_distance_0039 <= 874568;
    i_distance_0040 <= 583498;
    i_distance_0041 <= 362571;
    i_distance_0042 <= 1015499;
    i_distance_0043 <= 15700;
    i_distance_0044 <= 915540;
    i_distance_0045 <= 873430;
    i_distance_0046 <= 11991;
    i_distance_0047 <= 555610;
    i_distance_0048 <= 388826;
    i_distance_0049 <= 346330;
    i_distance_0050 <= 275423;
    i_distance_0051 <= 404320;
    i_distance_0052 <= 252898;
    i_distance_0053 <= 829795;
    i_distance_0054 <= 288615;
    i_distance_0055 <= 401000;
    i_distance_0056 <= 372073;
    i_distance_0057 <= 174702;
    i_distance_0058 <= 354287;
    i_distance_0059 <= 285552;
    i_distance_0060 <= 335349;
    i_distance_0061 <= 51574;
    i_distance_0062 <= 251768;
    i_distance_0063 <= 280191;
    correct_answer <= 11991;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 429184;
    i_distance_0001 <= 434945;
    i_distance_0002 <= 74375;
    i_distance_0003 <= 452615;
    i_distance_0004 <= 183949;
    i_distance_0005 <= 693393;
    i_distance_0006 <= 453012;
    i_distance_0007 <= 723221;
    i_distance_0008 <= 812182;
    i_distance_0009 <= 628892;
    i_distance_0010 <= 530077;
    i_distance_0011 <= 70049;
    i_distance_0012 <= 485921;
    i_distance_0013 <= 690595;
    i_distance_0014 <= 614438;
    i_distance_0015 <= 70695;
    i_distance_0016 <= 427559;
    i_distance_0017 <= 889513;
    i_distance_0018 <= 544169;
    i_distance_0019 <= 215851;
    i_distance_0020 <= 495150;
    i_distance_0021 <= 943791;
    i_distance_0022 <= 292145;
    i_distance_0023 <= 93490;
    i_distance_0024 <= 914738;
    i_distance_0025 <= 460852;
    i_distance_0026 <= 1035317;
    i_distance_0027 <= 860727;
    i_distance_0028 <= 836538;
    i_distance_0029 <= 390331;
    i_distance_0030 <= 774460;
    i_distance_0031 <= 1039805;
    i_distance_0032 <= 416958;
    i_distance_0033 <= 39486;
    i_distance_0034 <= 30139;
    i_distance_0035 <= 86463;
    i_distance_0036 <= 959426;
    i_distance_0037 <= 781762;
    i_distance_0038 <= 274491;
    i_distance_0039 <= 751559;
    i_distance_0040 <= 701390;
    i_distance_0041 <= 654926;
    i_distance_0042 <= 362451;
    i_distance_0043 <= 218964;
    i_distance_0044 <= 439765;
    i_distance_0045 <= 534355;
    i_distance_0046 <= 35289;
    i_distance_0047 <= 655194;
    i_distance_0048 <= 341338;
    i_distance_0049 <= 819703;
    i_distance_0050 <= 983653;
    i_distance_0051 <= 415462;
    i_distance_0052 <= 144997;
    i_distance_0053 <= 793446;
    i_distance_0054 <= 293227;
    i_distance_0055 <= 867054;
    i_distance_0056 <= 589294;
    i_distance_0057 <= 811248;
    i_distance_0058 <= 883697;
    i_distance_0059 <= 133495;
    i_distance_0060 <= 58232;
    i_distance_0061 <= 638201;
    i_distance_0062 <= 755707;
    i_distance_0063 <= 385020;
    correct_answer <= 30139;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 27778;
    i_distance_0001 <= 919172;
    i_distance_0002 <= 146309;
    i_distance_0003 <= 703494;
    i_distance_0004 <= 136456;
    i_distance_0005 <= 91147;
    i_distance_0006 <= 97036;
    i_distance_0007 <= 373389;
    i_distance_0008 <= 898830;
    i_distance_0009 <= 122639;
    i_distance_0010 <= 925585;
    i_distance_0011 <= 865041;
    i_distance_0012 <= 560787;
    i_distance_0013 <= 353683;
    i_distance_0014 <= 294553;
    i_distance_0015 <= 518812;
    i_distance_0016 <= 375197;
    i_distance_0017 <= 295838;
    i_distance_0018 <= 901795;
    i_distance_0019 <= 701604;
    i_distance_0020 <= 2595;
    i_distance_0021 <= 152361;
    i_distance_0022 <= 280617;
    i_distance_0023 <= 707884;
    i_distance_0024 <= 370734;
    i_distance_0025 <= 711343;
    i_distance_0026 <= 499760;
    i_distance_0027 <= 581681;
    i_distance_0028 <= 1035568;
    i_distance_0029 <= 639667;
    i_distance_0030 <= 165172;
    i_distance_0031 <= 492854;
    i_distance_0032 <= 586294;
    i_distance_0033 <= 478396;
    i_distance_0034 <= 901693;
    i_distance_0035 <= 764224;
    i_distance_0036 <= 563907;
    i_distance_0037 <= 201796;
    i_distance_0038 <= 797639;
    i_distance_0039 <= 558156;
    i_distance_0040 <= 923597;
    i_distance_0041 <= 191310;
    i_distance_0042 <= 35919;
    i_distance_0043 <= 783955;
    i_distance_0044 <= 306133;
    i_distance_0045 <= 497625;
    i_distance_0046 <= 103519;
    i_distance_0047 <= 570464;
    i_distance_0048 <= 713444;
    i_distance_0049 <= 259941;
    i_distance_0050 <= 780516;
    i_distance_0051 <= 793194;
    i_distance_0052 <= 204266;
    i_distance_0053 <= 113772;
    i_distance_0054 <= 892781;
    i_distance_0055 <= 194032;
    i_distance_0056 <= 475760;
    i_distance_0057 <= 136307;
    i_distance_0058 <= 49525;
    i_distance_0059 <= 5750;
    i_distance_0060 <= 659192;
    i_distance_0061 <= 71291;
    i_distance_0062 <= 702844;
    i_distance_0063 <= 921470;
    correct_answer <= 2595;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 170628;
    i_distance_0001 <= 109063;
    i_distance_0002 <= 246794;
    i_distance_0003 <= 535565;
    i_distance_0004 <= 796943;
    i_distance_0005 <= 350096;
    i_distance_0006 <= 513169;
    i_distance_0007 <= 462609;
    i_distance_0008 <= 178064;
    i_distance_0009 <= 499088;
    i_distance_0010 <= 323605;
    i_distance_0011 <= 198160;
    i_distance_0012 <= 945946;
    i_distance_0013 <= 854428;
    i_distance_0014 <= 541343;
    i_distance_0015 <= 686879;
    i_distance_0016 <= 222244;
    i_distance_0017 <= 790692;
    i_distance_0018 <= 771754;
    i_distance_0019 <= 888620;
    i_distance_0020 <= 938028;
    i_distance_0021 <= 613038;
    i_distance_0022 <= 672432;
    i_distance_0023 <= 1021496;
    i_distance_0024 <= 401593;
    i_distance_0025 <= 754234;
    i_distance_0026 <= 215610;
    i_distance_0027 <= 693309;
    i_distance_0028 <= 737086;
    i_distance_0029 <= 738493;
    i_distance_0030 <= 660034;
    i_distance_0031 <= 436803;
    i_distance_0032 <= 1035715;
    i_distance_0033 <= 782661;
    i_distance_0034 <= 810694;
    i_distance_0035 <= 984642;
    i_distance_0036 <= 805199;
    i_distance_0037 <= 670032;
    i_distance_0038 <= 215633;
    i_distance_0039 <= 115537;
    i_distance_0040 <= 490837;
    i_distance_0041 <= 467542;
    i_distance_0042 <= 71386;
    i_distance_0043 <= 610398;
    i_distance_0044 <= 538464;
    i_distance_0045 <= 678114;
    i_distance_0046 <= 585573;
    i_distance_0047 <= 996455;
    i_distance_0048 <= 137448;
    i_distance_0049 <= 62312;
    i_distance_0050 <= 1001962;
    i_distance_0051 <= 7787;
    i_distance_0052 <= 631403;
    i_distance_0053 <= 410601;
    i_distance_0054 <= 218730;
    i_distance_0055 <= 334831;
    i_distance_0056 <= 508015;
    i_distance_0057 <= 8433;
    i_distance_0058 <= 1021685;
    i_distance_0059 <= 172150;
    i_distance_0060 <= 939257;
    i_distance_0061 <= 984443;
    i_distance_0062 <= 797949;
    i_distance_0063 <= 603390;
    correct_answer <= 7787;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 422539;
    i_distance_0001 <= 286987;
    i_distance_0002 <= 110091;
    i_distance_0003 <= 1010958;
    i_distance_0004 <= 612619;
    i_distance_0005 <= 98064;
    i_distance_0006 <= 548880;
    i_distance_0007 <= 337298;
    i_distance_0008 <= 479379;
    i_distance_0009 <= 817938;
    i_distance_0010 <= 558606;
    i_distance_0011 <= 440464;
    i_distance_0012 <= 211607;
    i_distance_0013 <= 264090;
    i_distance_0014 <= 835355;
    i_distance_0015 <= 509596;
    i_distance_0016 <= 763685;
    i_distance_0017 <= 3110;
    i_distance_0018 <= 658602;
    i_distance_0019 <= 478638;
    i_distance_0020 <= 237233;
    i_distance_0021 <= 770868;
    i_distance_0022 <= 742708;
    i_distance_0023 <= 580790;
    i_distance_0024 <= 31159;
    i_distance_0025 <= 780286;
    i_distance_0026 <= 482107;
    i_distance_0027 <= 575676;
    i_distance_0028 <= 431549;
    i_distance_0029 <= 472380;
    i_distance_0030 <= 619711;
    i_distance_0031 <= 146624;
    i_distance_0032 <= 762689;
    i_distance_0033 <= 125376;
    i_distance_0034 <= 899136;
    i_distance_0035 <= 967876;
    i_distance_0036 <= 724163;
    i_distance_0037 <= 1035465;
    i_distance_0038 <= 493129;
    i_distance_0039 <= 58959;
    i_distance_0040 <= 809552;
    i_distance_0041 <= 339280;
    i_distance_0042 <= 549971;
    i_distance_0043 <= 585684;
    i_distance_0044 <= 1012566;
    i_distance_0045 <= 439774;
    i_distance_0046 <= 1003743;
    i_distance_0047 <= 516191;
    i_distance_0048 <= 166368;
    i_distance_0049 <= 577504;
    i_distance_0050 <= 893411;
    i_distance_0051 <= 542819;
    i_distance_0052 <= 288229;
    i_distance_0053 <= 573032;
    i_distance_0054 <= 690664;
    i_distance_0055 <= 353258;
    i_distance_0056 <= 988785;
    i_distance_0057 <= 89716;
    i_distance_0058 <= 944117;
    i_distance_0059 <= 75124;
    i_distance_0060 <= 613368;
    i_distance_0061 <= 814204;
    i_distance_0062 <= 588798;
    i_distance_0063 <= 1012991;
    correct_answer <= 3110;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 136064;
    i_distance_0001 <= 174850;
    i_distance_0002 <= 262915;
    i_distance_0003 <= 647171;
    i_distance_0004 <= 928389;
    i_distance_0005 <= 726787;
    i_distance_0006 <= 626819;
    i_distance_0007 <= 159369;
    i_distance_0008 <= 438028;
    i_distance_0009 <= 1019918;
    i_distance_0010 <= 179599;
    i_distance_0011 <= 592144;
    i_distance_0012 <= 17422;
    i_distance_0013 <= 1018772;
    i_distance_0014 <= 492820;
    i_distance_0015 <= 880792;
    i_distance_0016 <= 766619;
    i_distance_0017 <= 498460;
    i_distance_0018 <= 382244;
    i_distance_0019 <= 280357;
    i_distance_0020 <= 477861;
    i_distance_0021 <= 380968;
    i_distance_0022 <= 856616;
    i_distance_0023 <= 238891;
    i_distance_0024 <= 470572;
    i_distance_0025 <= 463024;
    i_distance_0026 <= 142769;
    i_distance_0027 <= 353713;
    i_distance_0028 <= 922163;
    i_distance_0029 <= 711092;
    i_distance_0030 <= 552502;
    i_distance_0031 <= 588214;
    i_distance_0032 <= 129210;
    i_distance_0033 <= 896061;
    i_distance_0034 <= 451005;
    i_distance_0035 <= 873405;
    i_distance_0036 <= 23870;
    i_distance_0037 <= 859464;
    i_distance_0038 <= 820937;
    i_distance_0039 <= 655563;
    i_distance_0040 <= 1022159;
    i_distance_0041 <= 684496;
    i_distance_0042 <= 766161;
    i_distance_0043 <= 511058;
    i_distance_0044 <= 587605;
    i_distance_0045 <= 326230;
    i_distance_0046 <= 1009238;
    i_distance_0047 <= 1044952;
    i_distance_0048 <= 255448;
    i_distance_0049 <= 1045338;
    i_distance_0050 <= 765054;
    i_distance_0051 <= 41052;
    i_distance_0052 <= 144606;
    i_distance_0053 <= 534111;
    i_distance_0054 <= 31456;
    i_distance_0055 <= 469986;
    i_distance_0056 <= 670575;
    i_distance_0057 <= 191344;
    i_distance_0058 <= 542706;
    i_distance_0059 <= 125170;
    i_distance_0060 <= 550261;
    i_distance_0061 <= 971511;
    i_distance_0062 <= 339194;
    i_distance_0063 <= 43390;
    correct_answer <= 17422;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 638080;
    i_distance_0001 <= 71041;
    i_distance_0002 <= 317313;
    i_distance_0003 <= 670211;
    i_distance_0004 <= 1033859;
    i_distance_0005 <= 292485;
    i_distance_0006 <= 800006;
    i_distance_0007 <= 1047172;
    i_distance_0008 <= 291209;
    i_distance_0009 <= 389260;
    i_distance_0010 <= 525581;
    i_distance_0011 <= 1026702;
    i_distance_0012 <= 328975;
    i_distance_0013 <= 944787;
    i_distance_0014 <= 250646;
    i_distance_0015 <= 231320;
    i_distance_0016 <= 14233;
    i_distance_0017 <= 227226;
    i_distance_0018 <= 317082;
    i_distance_0019 <= 968990;
    i_distance_0020 <= 335647;
    i_distance_0021 <= 163230;
    i_distance_0022 <= 558115;
    i_distance_0023 <= 1020580;
    i_distance_0024 <= 635174;
    i_distance_0025 <= 64687;
    i_distance_0026 <= 963121;
    i_distance_0027 <= 766644;
    i_distance_0028 <= 740405;
    i_distance_0029 <= 1029687;
    i_distance_0030 <= 746936;
    i_distance_0031 <= 125628;
    i_distance_0032 <= 226877;
    i_distance_0033 <= 1000770;
    i_distance_0034 <= 698698;
    i_distance_0035 <= 690507;
    i_distance_0036 <= 20812;
    i_distance_0037 <= 997580;
    i_distance_0038 <= 1039179;
    i_distance_0039 <= 458832;
    i_distance_0040 <= 983506;
    i_distance_0041 <= 230099;
    i_distance_0042 <= 678227;
    i_distance_0043 <= 940757;
    i_distance_0044 <= 377686;
    i_distance_0045 <= 863575;
    i_distance_0046 <= 714845;
    i_distance_0047 <= 569182;
    i_distance_0048 <= 978141;
    i_distance_0049 <= 430817;
    i_distance_0050 <= 230242;
    i_distance_0051 <= 191073;
    i_distance_0052 <= 218470;
    i_distance_0053 <= 1039846;
    i_distance_0054 <= 833775;
    i_distance_0055 <= 338415;
    i_distance_0056 <= 266097;
    i_distance_0057 <= 612596;
    i_distance_0058 <= 28407;
    i_distance_0059 <= 102776;
    i_distance_0060 <= 633;
    i_distance_0061 <= 928635;
    i_distance_0062 <= 852989;
    i_distance_0063 <= 970751;
    correct_answer <= 633;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 660356;
    i_distance_0001 <= 341387;
    i_distance_0002 <= 815116;
    i_distance_0003 <= 1004427;
    i_distance_0004 <= 522388;
    i_distance_0005 <= 735893;
    i_distance_0006 <= 787605;
    i_distance_0007 <= 864920;
    i_distance_0008 <= 481695;
    i_distance_0009 <= 595871;
    i_distance_0010 <= 782113;
    i_distance_0011 <= 784674;
    i_distance_0012 <= 148128;
    i_distance_0013 <= 133670;
    i_distance_0014 <= 265639;
    i_distance_0015 <= 261672;
    i_distance_0016 <= 431785;
    i_distance_0017 <= 404010;
    i_distance_0018 <= 745003;
    i_distance_0019 <= 908204;
    i_distance_0020 <= 898350;
    i_distance_0021 <= 594351;
    i_distance_0022 <= 81455;
    i_distance_0023 <= 634160;
    i_distance_0024 <= 743857;
    i_distance_0025 <= 127157;
    i_distance_0026 <= 489531;
    i_distance_0027 <= 693436;
    i_distance_0028 <= 122173;
    i_distance_0029 <= 540992;
    i_distance_0030 <= 731968;
    i_distance_0031 <= 61635;
    i_distance_0032 <= 570053;
    i_distance_0033 <= 25670;
    i_distance_0034 <= 994119;
    i_distance_0035 <= 287558;
    i_distance_0036 <= 467657;
    i_distance_0037 <= 564813;
    i_distance_0038 <= 851918;
    i_distance_0039 <= 367868;
    i_distance_0040 <= 746198;
    i_distance_0041 <= 549078;
    i_distance_0042 <= 548182;
    i_distance_0043 <= 720217;
    i_distance_0044 <= 209242;
    i_distance_0045 <= 730840;
    i_distance_0046 <= 74080;
    i_distance_0047 <= 187745;
    i_distance_0048 <= 741347;
    i_distance_0049 <= 1028580;
    i_distance_0050 <= 81124;
    i_distance_0051 <= 659940;
    i_distance_0052 <= 521828;
    i_distance_0053 <= 1030247;
    i_distance_0054 <= 1006570;
    i_distance_0055 <= 539755;
    i_distance_0056 <= 450288;
    i_distance_0057 <= 738801;
    i_distance_0058 <= 666101;
    i_distance_0059 <= 23414;
    i_distance_0060 <= 77943;
    i_distance_0061 <= 372091;
    i_distance_0062 <= 346620;
    i_distance_0063 <= 417279;
    correct_answer <= 23414;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 642567;
    i_distance_0001 <= 887815;
    i_distance_0002 <= 260234;
    i_distance_0003 <= 744844;
    i_distance_0004 <= 299021;
    i_distance_0005 <= 710541;
    i_distance_0006 <= 745873;
    i_distance_0007 <= 1170;
    i_distance_0008 <= 526995;
    i_distance_0009 <= 267414;
    i_distance_0010 <= 528151;
    i_distance_0011 <= 485656;
    i_distance_0012 <= 474009;
    i_distance_0013 <= 38808;
    i_distance_0014 <= 11671;
    i_distance_0015 <= 367772;
    i_distance_0016 <= 658462;
    i_distance_0017 <= 154142;
    i_distance_0018 <= 63648;
    i_distance_0019 <= 808993;
    i_distance_0020 <= 49056;
    i_distance_0021 <= 12318;
    i_distance_0022 <= 626855;
    i_distance_0023 <= 798119;
    i_distance_0024 <= 518696;
    i_distance_0025 <= 580139;
    i_distance_0026 <= 1024556;
    i_distance_0027 <= 103723;
    i_distance_0028 <= 359089;
    i_distance_0029 <= 769591;
    i_distance_0030 <= 237756;
    i_distance_0031 <= 556989;
    i_distance_0032 <= 105929;
    i_distance_0033 <= 840010;
    i_distance_0034 <= 649034;
    i_distance_0035 <= 253644;
    i_distance_0036 <= 747977;
    i_distance_0037 <= 704212;
    i_distance_0038 <= 1031381;
    i_distance_0039 <= 323029;
    i_distance_0040 <= 571863;
    i_distance_0041 <= 368728;
    i_distance_0042 <= 842199;
    i_distance_0043 <= 577245;
    i_distance_0044 <= 181086;
    i_distance_0045 <= 564958;
    i_distance_0046 <= 141283;
    i_distance_0047 <= 665956;
    i_distance_0048 <= 64741;
    i_distance_0049 <= 472934;
    i_distance_0050 <= 835811;
    i_distance_0051 <= 338532;
    i_distance_0052 <= 728303;
    i_distance_0053 <= 353392;
    i_distance_0054 <= 999025;
    i_distance_0055 <= 1008370;
    i_distance_0056 <= 416370;
    i_distance_0057 <= 90609;
    i_distance_0058 <= 742261;
    i_distance_0059 <= 219123;
    i_distance_0060 <= 102904;
    i_distance_0061 <= 845305;
    i_distance_0062 <= 784252;
    i_distance_0063 <= 165503;
    correct_answer <= 1170;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 47616;
    i_distance_0001 <= 862209;
    i_distance_0002 <= 430979;
    i_distance_0003 <= 320004;
    i_distance_0004 <= 459397;
    i_distance_0005 <= 207747;
    i_distance_0006 <= 894860;
    i_distance_0007 <= 397326;
    i_distance_0008 <= 243983;
    i_distance_0009 <= 663441;
    i_distance_0010 <= 173970;
    i_distance_0011 <= 984081;
    i_distance_0012 <= 745365;
    i_distance_0013 <= 104090;
    i_distance_0014 <= 620575;
    i_distance_0015 <= 154276;
    i_distance_0016 <= 546340;
    i_distance_0017 <= 943656;
    i_distance_0018 <= 1022121;
    i_distance_0019 <= 941999;
    i_distance_0020 <= 419123;
    i_distance_0021 <= 213558;
    i_distance_0022 <= 739513;
    i_distance_0023 <= 936511;
    i_distance_0024 <= 513984;
    i_distance_0025 <= 868929;
    i_distance_0026 <= 183106;
    i_distance_0027 <= 465091;
    i_distance_0028 <= 176833;
    i_distance_0029 <= 249797;
    i_distance_0030 <= 390472;
    i_distance_0031 <= 132425;
    i_distance_0032 <= 816968;
    i_distance_0033 <= 68043;
    i_distance_0034 <= 1031756;
    i_distance_0035 <= 622669;
    i_distance_0036 <= 79054;
    i_distance_0037 <= 355705;
    i_distance_0038 <= 272848;
    i_distance_0039 <= 107216;
    i_distance_0040 <= 161874;
    i_distance_0041 <= 437195;
    i_distance_0042 <= 735700;
    i_distance_0043 <= 122711;
    i_distance_0044 <= 61278;
    i_distance_0045 <= 489060;
    i_distance_0046 <= 71652;
    i_distance_0047 <= 351204;
    i_distance_0048 <= 844775;
    i_distance_0049 <= 993511;
    i_distance_0050 <= 284905;
    i_distance_0051 <= 26474;
    i_distance_0052 <= 116966;
    i_distance_0053 <= 672748;
    i_distance_0054 <= 225380;
    i_distance_0055 <= 446190;
    i_distance_0056 <= 411755;
    i_distance_0057 <= 174062;
    i_distance_0058 <= 520562;
    i_distance_0059 <= 122227;
    i_distance_0060 <= 755186;
    i_distance_0061 <= 814712;
    i_distance_0062 <= 537465;
    i_distance_0063 <= 14586;
    correct_answer <= 14586;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 667136;
    i_distance_0001 <= 736257;
    i_distance_0002 <= 773377;
    i_distance_0003 <= 358785;
    i_distance_0004 <= 960257;
    i_distance_0005 <= 945416;
    i_distance_0006 <= 68876;
    i_distance_0007 <= 913678;
    i_distance_0008 <= 79502;
    i_distance_0009 <= 952056;
    i_distance_0010 <= 626319;
    i_distance_0011 <= 805012;
    i_distance_0012 <= 1047190;
    i_distance_0013 <= 939928;
    i_distance_0014 <= 171036;
    i_distance_0015 <= 330910;
    i_distance_0016 <= 788129;
    i_distance_0017 <= 585634;
    i_distance_0018 <= 715813;
    i_distance_0019 <= 732454;
    i_distance_0020 <= 316837;
    i_distance_0021 <= 674086;
    i_distance_0022 <= 108971;
    i_distance_0023 <= 139693;
    i_distance_0024 <= 897967;
    i_distance_0025 <= 376880;
    i_distance_0026 <= 578992;
    i_distance_0027 <= 338226;
    i_distance_0028 <= 433586;
    i_distance_0029 <= 448308;
    i_distance_0030 <= 662197;
    i_distance_0031 <= 515760;
    i_distance_0032 <= 406584;
    i_distance_0033 <= 247737;
    i_distance_0034 <= 710968;
    i_distance_0035 <= 400187;
    i_distance_0036 <= 900285;
    i_distance_0037 <= 94013;
    i_distance_0038 <= 680513;
    i_distance_0039 <= 688579;
    i_distance_0040 <= 354632;
    i_distance_0041 <= 351185;
    i_distance_0042 <= 317397;
    i_distance_0043 <= 905429;
    i_distance_0044 <= 130903;
    i_distance_0045 <= 750425;
    i_distance_0046 <= 229854;
    i_distance_0047 <= 231395;
    i_distance_0048 <= 39396;
    i_distance_0049 <= 701283;
    i_distance_0050 <= 171110;
    i_distance_0051 <= 9960;
    i_distance_0052 <= 265961;
    i_distance_0053 <= 892138;
    i_distance_0054 <= 516331;
    i_distance_0055 <= 494828;
    i_distance_0056 <= 105321;
    i_distance_0057 <= 95983;
    i_distance_0058 <= 437489;
    i_distance_0059 <= 461555;
    i_distance_0060 <= 18550;
    i_distance_0061 <= 521591;
    i_distance_0062 <= 51704;
    i_distance_0063 <= 358271;
    correct_answer <= 9960;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 615168;
    i_distance_0001 <= 58754;
    i_distance_0002 <= 408197;
    i_distance_0003 <= 376837;
    i_distance_0004 <= 224010;
    i_distance_0005 <= 255372;
    i_distance_0006 <= 1023501;
    i_distance_0007 <= 218124;
    i_distance_0008 <= 389394;
    i_distance_0009 <= 337555;
    i_distance_0010 <= 507925;
    i_distance_0011 <= 486294;
    i_distance_0012 <= 26389;
    i_distance_0013 <= 729368;
    i_distance_0014 <= 878745;
    i_distance_0015 <= 439199;
    i_distance_0016 <= 920992;
    i_distance_0017 <= 310948;
    i_distance_0018 <= 158373;
    i_distance_0019 <= 231078;
    i_distance_0020 <= 676264;
    i_distance_0021 <= 11944;
    i_distance_0022 <= 951978;
    i_distance_0023 <= 63403;
    i_distance_0024 <= 480942;
    i_distance_0025 <= 734895;
    i_distance_0026 <= 220976;
    i_distance_0027 <= 745137;
    i_distance_0028 <= 1716;
    i_distance_0029 <= 877366;
    i_distance_0030 <= 179896;
    i_distance_0031 <= 662458;
    i_distance_0032 <= 872507;
    i_distance_0033 <= 915134;
    i_distance_0034 <= 387137;
    i_distance_0035 <= 68034;
    i_distance_0036 <= 558532;
    i_distance_0037 <= 81733;
    i_distance_0038 <= 147654;
    i_distance_0039 <= 159303;
    i_distance_0040 <= 794057;
    i_distance_0041 <= 1044684;
    i_distance_0042 <= 843853;
    i_distance_0043 <= 589646;
    i_distance_0044 <= 841679;
    i_distance_0045 <= 760273;
    i_distance_0046 <= 686547;
    i_distance_0047 <= 741336;
    i_distance_0048 <= 964825;
    i_distance_0049 <= 709593;
    i_distance_0050 <= 796768;
    i_distance_0051 <= 65761;
    i_distance_0052 <= 402405;
    i_distance_0053 <= 716389;
    i_distance_0054 <= 281701;
    i_distance_0055 <= 15464;
    i_distance_0056 <= 635881;
    i_distance_0057 <= 709996;
    i_distance_0058 <= 243952;
    i_distance_0059 <= 803826;
    i_distance_0060 <= 308089;
    i_distance_0061 <= 1032698;
    i_distance_0062 <= 543484;
    i_distance_0063 <= 972029;
    correct_answer <= 1716;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 729088;
    i_distance_0001 <= 698370;
    i_distance_0002 <= 99075;
    i_distance_0003 <= 828548;
    i_distance_0004 <= 681991;
    i_distance_0005 <= 579082;
    i_distance_0006 <= 569612;
    i_distance_0007 <= 717967;
    i_distance_0008 <= 460821;
    i_distance_0009 <= 274583;
    i_distance_0010 <= 261400;
    i_distance_0011 <= 574363;
    i_distance_0012 <= 328732;
    i_distance_0013 <= 454685;
    i_distance_0014 <= 652317;
    i_distance_0015 <= 822815;
    i_distance_0016 <= 927520;
    i_distance_0017 <= 409248;
    i_distance_0018 <= 520738;
    i_distance_0019 <= 729377;
    i_distance_0020 <= 371238;
    i_distance_0021 <= 761769;
    i_distance_0022 <= 152877;
    i_distance_0023 <= 1021743;
    i_distance_0024 <= 841781;
    i_distance_0025 <= 110518;
    i_distance_0026 <= 940597;
    i_distance_0027 <= 143800;
    i_distance_0028 <= 587701;
    i_distance_0029 <= 903738;
    i_distance_0030 <= 108219;
    i_distance_0031 <= 981565;
    i_distance_0032 <= 969535;
    i_distance_0033 <= 383612;
    i_distance_0034 <= 272449;
    i_distance_0035 <= 962499;
    i_distance_0036 <= 34502;
    i_distance_0037 <= 967112;
    i_distance_0038 <= 357067;
    i_distance_0039 <= 884300;
    i_distance_0040 <= 466253;
    i_distance_0041 <= 728013;
    i_distance_0042 <= 910284;
    i_distance_0043 <= 61003;
    i_distance_0044 <= 16977;
    i_distance_0045 <= 862164;
    i_distance_0046 <= 980438;
    i_distance_0047 <= 396761;
    i_distance_0048 <= 444634;
    i_distance_0049 <= 682329;
    i_distance_0050 <= 246620;
    i_distance_0051 <= 237918;
    i_distance_0052 <= 756706;
    i_distance_0053 <= 389859;
    i_distance_0054 <= 912226;
    i_distance_0055 <= 383079;
    i_distance_0056 <= 801900;
    i_distance_0057 <= 381165;
    i_distance_0058 <= 388462;
    i_distance_0059 <= 1015152;
    i_distance_0060 <= 533236;
    i_distance_0061 <= 949369;
    i_distance_0062 <= 914684;
    i_distance_0063 <= 310143;
    correct_answer <= 16977;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 52225;
    i_distance_0001 <= 386309;
    i_distance_0002 <= 1033349;
    i_distance_0003 <= 758277;
    i_distance_0004 <= 336648;
    i_distance_0005 <= 960011;
    i_distance_0006 <= 850188;
    i_distance_0007 <= 445075;
    i_distance_0008 <= 887571;
    i_distance_0009 <= 956952;
    i_distance_0010 <= 872089;
    i_distance_0011 <= 600347;
    i_distance_0012 <= 557981;
    i_distance_0013 <= 303645;
    i_distance_0014 <= 598943;
    i_distance_0015 <= 768376;
    i_distance_0016 <= 347301;
    i_distance_0017 <= 416677;
    i_distance_0018 <= 47142;
    i_distance_0019 <= 101290;
    i_distance_0020 <= 823212;
    i_distance_0021 <= 918449;
    i_distance_0022 <= 141106;
    i_distance_0023 <= 796211;
    i_distance_0024 <= 702644;
    i_distance_0025 <= 650164;
    i_distance_0026 <= 1024561;
    i_distance_0027 <= 127539;
    i_distance_0028 <= 56372;
    i_distance_0029 <= 169787;
    i_distance_0030 <= 742846;
    i_distance_0031 <= 437827;
    i_distance_0032 <= 997830;
    i_distance_0033 <= 228423;
    i_distance_0034 <= 27081;
    i_distance_0035 <= 1024713;
    i_distance_0036 <= 482765;
    i_distance_0037 <= 680145;
    i_distance_0038 <= 562258;
    i_distance_0039 <= 967507;
    i_distance_0040 <= 111700;
    i_distance_0041 <= 253908;
    i_distance_0042 <= 513367;
    i_distance_0043 <= 352346;
    i_distance_0044 <= 611674;
    i_distance_0045 <= 762337;
    i_distance_0046 <= 389218;
    i_distance_0047 <= 100835;
    i_distance_0048 <= 1008355;
    i_distance_0049 <= 529509;
    i_distance_0050 <= 395366;
    i_distance_0051 <= 293988;
    i_distance_0052 <= 154089;
    i_distance_0053 <= 907370;
    i_distance_0054 <= 320618;
    i_distance_0055 <= 937708;
    i_distance_0056 <= 970221;
    i_distance_0057 <= 45684;
    i_distance_0058 <= 149109;
    i_distance_0059 <= 920565;
    i_distance_0060 <= 728568;
    i_distance_0061 <= 1018361;
    i_distance_0062 <= 190077;
    i_distance_0063 <= 688639;
    correct_answer <= 27081;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 840577;
    i_distance_0001 <= 63234;
    i_distance_0002 <= 965249;
    i_distance_0003 <= 430852;
    i_distance_0004 <= 630151;
    i_distance_0005 <= 136073;
    i_distance_0006 <= 268554;
    i_distance_0007 <= 955657;
    i_distance_0008 <= 900748;
    i_distance_0009 <= 643468;
    i_distance_0010 <= 939531;
    i_distance_0011 <= 160273;
    i_distance_0012 <= 256915;
    i_distance_0013 <= 286101;
    i_distance_0014 <= 224281;
    i_distance_0015 <= 441247;
    i_distance_0016 <= 7839;
    i_distance_0017 <= 231073;
    i_distance_0018 <= 928673;
    i_distance_0019 <= 1038884;
    i_distance_0020 <= 480425;
    i_distance_0021 <= 803881;
    i_distance_0022 <= 190125;
    i_distance_0023 <= 614195;
    i_distance_0024 <= 914228;
    i_distance_0025 <= 430902;
    i_distance_0026 <= 98103;
    i_distance_0027 <= 408632;
    i_distance_0028 <= 1038905;
    i_distance_0029 <= 772281;
    i_distance_0030 <= 343867;
    i_distance_0031 <= 956475;
    i_distance_0032 <= 770493;
    i_distance_0033 <= 11710;
    i_distance_0034 <= 356031;
    i_distance_0035 <= 552262;
    i_distance_0036 <= 655949;
    i_distance_0037 <= 814286;
    i_distance_0038 <= 530614;
    i_distance_0039 <= 3548;
    i_distance_0040 <= 159452;
    i_distance_0041 <= 501341;
    i_distance_0042 <= 841823;
    i_distance_0043 <= 68704;
    i_distance_0044 <= 136286;
    i_distance_0045 <= 571232;
    i_distance_0046 <= 412086;
    i_distance_0047 <= 691297;
    i_distance_0048 <= 837221;
    i_distance_0049 <= 559077;
    i_distance_0050 <= 247781;
    i_distance_0051 <= 816360;
    i_distance_0052 <= 110440;
    i_distance_0053 <= 757610;
    i_distance_0054 <= 468202;
    i_distance_0055 <= 42733;
    i_distance_0056 <= 500846;
    i_distance_0057 <= 530159;
    i_distance_0058 <= 152945;
    i_distance_0059 <= 122738;
    i_distance_0060 <= 90355;
    i_distance_0061 <= 536690;
    i_distance_0062 <= 605817;
    i_distance_0063 <= 743807;
    correct_answer <= 3548;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 122372;
    i_distance_0001 <= 1029764;
    i_distance_0002 <= 281478;
    i_distance_0003 <= 230532;
    i_distance_0004 <= 208008;
    i_distance_0005 <= 399624;
    i_distance_0006 <= 817668;
    i_distance_0007 <= 12942;
    i_distance_0008 <= 875919;
    i_distance_0009 <= 987408;
    i_distance_0010 <= 345620;
    i_distance_0011 <= 799639;
    i_distance_0012 <= 373016;
    i_distance_0013 <= 746007;
    i_distance_0014 <= 35741;
    i_distance_0015 <= 805917;
    i_distance_0016 <= 780189;
    i_distance_0017 <= 894368;
    i_distance_0018 <= 17698;
    i_distance_0019 <= 243238;
    i_distance_0020 <= 1003942;
    i_distance_0021 <= 805164;
    i_distance_0022 <= 676396;
    i_distance_0023 <= 72492;
    i_distance_0024 <= 430133;
    i_distance_0025 <= 979766;
    i_distance_0026 <= 699831;
    i_distance_0027 <= 215740;
    i_distance_0028 <= 1000124;
    i_distance_0029 <= 213822;
    i_distance_0030 <= 153021;
    i_distance_0031 <= 987453;
    i_distance_0032 <= 708540;
    i_distance_0033 <= 623938;
    i_distance_0034 <= 977092;
    i_distance_0035 <= 389829;
    i_distance_0036 <= 1037381;
    i_distance_0037 <= 613960;
    i_distance_0038 <= 749129;
    i_distance_0039 <= 23372;
    i_distance_0040 <= 172109;
    i_distance_0041 <= 387151;
    i_distance_0042 <= 9168;
    i_distance_0043 <= 402386;
    i_distance_0044 <= 130259;
    i_distance_0045 <= 556244;
    i_distance_0046 <= 904152;
    i_distance_0047 <= 563299;
    i_distance_0048 <= 146660;
    i_distance_0049 <= 424423;
    i_distance_0050 <= 551656;
    i_distance_0051 <= 613097;
    i_distance_0052 <= 142698;
    i_distance_0053 <= 783594;
    i_distance_0054 <= 1043687;
    i_distance_0055 <= 114413;
    i_distance_0056 <= 253439;
    i_distance_0057 <= 780656;
    i_distance_0058 <= 417520;
    i_distance_0059 <= 609906;
    i_distance_0060 <= 931184;
    i_distance_0061 <= 500981;
    i_distance_0062 <= 353782;
    i_distance_0063 <= 494079;
    correct_answer <= 9168;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 527360;
    i_distance_0001 <= 513025;
    i_distance_0002 <= 976770;
    i_distance_0003 <= 566148;
    i_distance_0004 <= 236934;
    i_distance_0005 <= 146312;
    i_distance_0006 <= 97163;
    i_distance_0007 <= 1019916;
    i_distance_0008 <= 177934;
    i_distance_0009 <= 343825;
    i_distance_0010 <= 619411;
    i_distance_0011 <= 283391;
    i_distance_0012 <= 480534;
    i_distance_0013 <= 998295;
    i_distance_0014 <= 42518;
    i_distance_0015 <= 242589;
    i_distance_0016 <= 576288;
    i_distance_0017 <= 350625;
    i_distance_0018 <= 712355;
    i_distance_0019 <= 262179;
    i_distance_0020 <= 441893;
    i_distance_0021 <= 470056;
    i_distance_0022 <= 1022505;
    i_distance_0023 <= 705833;
    i_distance_0024 <= 366251;
    i_distance_0025 <= 531761;
    i_distance_0026 <= 260402;
    i_distance_0027 <= 346931;
    i_distance_0028 <= 332086;
    i_distance_0029 <= 883383;
    i_distance_0030 <= 389302;
    i_distance_0031 <= 508345;
    i_distance_0032 <= 216762;
    i_distance_0033 <= 1002743;
    i_distance_0034 <= 911614;
    i_distance_0035 <= 829634;
    i_distance_0036 <= 490436;
    i_distance_0037 <= 957637;
    i_distance_0038 <= 319176;
    i_distance_0039 <= 39624;
    i_distance_0040 <= 352840;
    i_distance_0041 <= 951243;
    i_distance_0042 <= 584523;
    i_distance_0043 <= 45771;
    i_distance_0044 <= 323278;
    i_distance_0045 <= 543487;
    i_distance_0046 <= 416599;
    i_distance_0047 <= 92376;
    i_distance_0048 <= 191963;
    i_distance_0049 <= 598876;
    i_distance_0050 <= 584668;
    i_distance_0051 <= 645212;
    i_distance_0052 <= 263521;
    i_distance_0053 <= 996452;
    i_distance_0054 <= 189416;
    i_distance_0055 <= 587761;
    i_distance_0056 <= 205170;
    i_distance_0057 <= 438514;
    i_distance_0058 <= 544628;
    i_distance_0059 <= 693878;
    i_distance_0060 <= 718199;
    i_distance_0061 <= 538492;
    i_distance_0062 <= 113662;
    i_distance_0063 <= 708095;
    correct_answer <= 39624;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 651269;
    i_distance_0001 <= 780678;
    i_distance_0002 <= 1047177;
    i_distance_0003 <= 863882;
    i_distance_0004 <= 453641;
    i_distance_0005 <= 302476;
    i_distance_0006 <= 213774;
    i_distance_0007 <= 528656;
    i_distance_0008 <= 74769;
    i_distance_0009 <= 344336;
    i_distance_0010 <= 670226;
    i_distance_0011 <= 817556;
    i_distance_0012 <= 1035920;
    i_distance_0013 <= 963990;
    i_distance_0014 <= 252436;
    i_distance_0015 <= 227347;
    i_distance_0016 <= 538263;
    i_distance_0017 <= 409370;
    i_distance_0018 <= 174110;
    i_distance_0019 <= 776478;
    i_distance_0020 <= 988702;
    i_distance_0021 <= 616136;
    i_distance_0022 <= 953508;
    i_distance_0023 <= 169126;
    i_distance_0024 <= 956070;
    i_distance_0025 <= 169896;
    i_distance_0026 <= 330153;
    i_distance_0027 <= 781225;
    i_distance_0028 <= 324781;
    i_distance_0029 <= 1005872;
    i_distance_0030 <= 459446;
    i_distance_0031 <= 164662;
    i_distance_0032 <= 400572;
    i_distance_0033 <= 720195;
    i_distance_0034 <= 979012;
    i_distance_0035 <= 378053;
    i_distance_0036 <= 8518;
    i_distance_0037 <= 776519;
    i_distance_0038 <= 867399;
    i_distance_0039 <= 916681;
    i_distance_0040 <= 714698;
    i_distance_0041 <= 58058;
    i_distance_0042 <= 212810;
    i_distance_0043 <= 586692;
    i_distance_0044 <= 737486;
    i_distance_0045 <= 279887;
    i_distance_0046 <= 331343;
    i_distance_0047 <= 660432;
    i_distance_0048 <= 120916;
    i_distance_0049 <= 878807;
    i_distance_0050 <= 965595;
    i_distance_0051 <= 637661;
    i_distance_0052 <= 132189;
    i_distance_0053 <= 1044319;
    i_distance_0054 <= 2525;
    i_distance_0055 <= 129634;
    i_distance_0056 <= 681575;
    i_distance_0057 <= 830568;
    i_distance_0058 <= 595306;
    i_distance_0059 <= 461679;
    i_distance_0060 <= 1009266;
    i_distance_0061 <= 327933;
    i_distance_0062 <= 267006;
    i_distance_0063 <= 462079;
    correct_answer <= 2525;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 688896;
    i_distance_0001 <= 974084;
    i_distance_0002 <= 481668;
    i_distance_0003 <= 989319;
    i_distance_0004 <= 250631;
    i_distance_0005 <= 136713;
    i_distance_0006 <= 713997;
    i_distance_0007 <= 224142;
    i_distance_0008 <= 731791;
    i_distance_0009 <= 681361;
    i_distance_0010 <= 272785;
    i_distance_0011 <= 426006;
    i_distance_0012 <= 439831;
    i_distance_0013 <= 581527;
    i_distance_0014 <= 413208;
    i_distance_0015 <= 630425;
    i_distance_0016 <= 564507;
    i_distance_0017 <= 176668;
    i_distance_0018 <= 998939;
    i_distance_0019 <= 958880;
    i_distance_0020 <= 900258;
    i_distance_0021 <= 874275;
    i_distance_0022 <= 989433;
    i_distance_0023 <= 498982;
    i_distance_0024 <= 366375;
    i_distance_0025 <= 783144;
    i_distance_0026 <= 868524;
    i_distance_0027 <= 654638;
    i_distance_0028 <= 242991;
    i_distance_0029 <= 107695;
    i_distance_0030 <= 966321;
    i_distance_0031 <= 169391;
    i_distance_0032 <= 454451;
    i_distance_0033 <= 330930;
    i_distance_0034 <= 789042;
    i_distance_0035 <= 546999;
    i_distance_0036 <= 376896;
    i_distance_0037 <= 579009;
    i_distance_0038 <= 65218;
    i_distance_0039 <= 813379;
    i_distance_0040 <= 17090;
    i_distance_0041 <= 1031417;
    i_distance_0042 <= 68672;
    i_distance_0043 <= 77000;
    i_distance_0044 <= 1019338;
    i_distance_0045 <= 250190;
    i_distance_0046 <= 615250;
    i_distance_0047 <= 325976;
    i_distance_0048 <= 40825;
    i_distance_0049 <= 888026;
    i_distance_0050 <= 845785;
    i_distance_0051 <= 185949;
    i_distance_0052 <= 674526;
    i_distance_0053 <= 619106;
    i_distance_0054 <= 364260;
    i_distance_0055 <= 834534;
    i_distance_0056 <= 250473;
    i_distance_0057 <= 666732;
    i_distance_0058 <= 332656;
    i_distance_0059 <= 469878;
    i_distance_0060 <= 465270;
    i_distance_0061 <= 983672;
    i_distance_0062 <= 204153;
    i_distance_0063 <= 508671;
    correct_answer <= 17090;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 201976;
    i_distance_0001 <= 69762;
    i_distance_0002 <= 551299;
    i_distance_0003 <= 695301;
    i_distance_0004 <= 957960;
    i_distance_0005 <= 382986;
    i_distance_0006 <= 1039246;
    i_distance_0007 <= 1023888;
    i_distance_0008 <= 894865;
    i_distance_0009 <= 1019411;
    i_distance_0010 <= 885779;
    i_distance_0011 <= 909718;
    i_distance_0012 <= 977559;
    i_distance_0013 <= 823575;
    i_distance_0014 <= 487582;
    i_distance_0015 <= 790560;
    i_distance_0016 <= 860195;
    i_distance_0017 <= 677796;
    i_distance_0018 <= 599334;
    i_distance_0019 <= 509095;
    i_distance_0020 <= 435114;
    i_distance_0021 <= 873130;
    i_distance_0022 <= 709548;
    i_distance_0023 <= 942767;
    i_distance_0024 <= 272562;
    i_distance_0025 <= 783794;
    i_distance_0026 <= 933688;
    i_distance_0027 <= 486205;
    i_distance_0028 <= 464961;
    i_distance_0029 <= 624452;
    i_distance_0030 <= 1016645;
    i_distance_0031 <= 468420;
    i_distance_0032 <= 873159;
    i_distance_0033 <= 112071;
    i_distance_0034 <= 747724;
    i_distance_0035 <= 495949;
    i_distance_0036 <= 917964;
    i_distance_0037 <= 720716;
    i_distance_0038 <= 807117;
    i_distance_0039 <= 278222;
    i_distance_0040 <= 464973;
    i_distance_0041 <= 647507;
    i_distance_0042 <= 88399;
    i_distance_0043 <= 794706;
    i_distance_0044 <= 6226;
    i_distance_0045 <= 850394;
    i_distance_0046 <= 848091;
    i_distance_0047 <= 1002077;
    i_distance_0048 <= 46814;
    i_distance_0049 <= 297313;
    i_distance_0050 <= 760419;
    i_distance_0051 <= 272740;
    i_distance_0052 <= 987493;
    i_distance_0053 <= 319848;
    i_distance_0054 <= 2793;
    i_distance_0055 <= 570987;
    i_distance_0056 <= 265582;
    i_distance_0057 <= 629999;
    i_distance_0058 <= 122993;
    i_distance_0059 <= 582131;
    i_distance_0060 <= 136437;
    i_distance_0061 <= 260728;
    i_distance_0062 <= 311673;
    i_distance_0063 <= 741242;
    correct_answer <= 2793;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 242689;
    i_distance_0001 <= 792194;
    i_distance_0002 <= 94338;
    i_distance_0003 <= 192642;
    i_distance_0004 <= 978692;
    i_distance_0005 <= 20614;
    i_distance_0006 <= 231811;
    i_distance_0007 <= 414341;
    i_distance_0008 <= 286209;
    i_distance_0009 <= 97934;
    i_distance_0010 <= 79503;
    i_distance_0011 <= 511889;
    i_distance_0012 <= 314003;
    i_distance_0013 <= 1016729;
    i_distance_0014 <= 744986;
    i_distance_0015 <= 221725;
    i_distance_0016 <= 769953;
    i_distance_0017 <= 157602;
    i_distance_0018 <= 657570;
    i_distance_0019 <= 825890;
    i_distance_0020 <= 767791;
    i_distance_0021 <= 245682;
    i_distance_0022 <= 294322;
    i_distance_0023 <= 862005;
    i_distance_0024 <= 866615;
    i_distance_0025 <= 113335;
    i_distance_0026 <= 69311;
    i_distance_0027 <= 592448;
    i_distance_0028 <= 37441;
    i_distance_0029 <= 617413;
    i_distance_0030 <= 332102;
    i_distance_0031 <= 371912;
    i_distance_0032 <= 966988;
    i_distance_0033 <= 654797;
    i_distance_0034 <= 185167;
    i_distance_0035 <= 785744;
    i_distance_0036 <= 90833;
    i_distance_0037 <= 809427;
    i_distance_0038 <= 116307;
    i_distance_0039 <= 149588;
    i_distance_0040 <= 1027030;
    i_distance_0041 <= 184151;
    i_distance_0042 <= 309079;
    i_distance_0043 <= 568408;
    i_distance_0044 <= 429779;
    i_distance_0045 <= 56917;
    i_distance_0046 <= 719315;
    i_distance_0047 <= 780125;
    i_distance_0048 <= 413816;
    i_distance_0049 <= 509025;
    i_distance_0050 <= 13410;
    i_distance_0051 <= 966503;
    i_distance_0052 <= 844007;
    i_distance_0053 <= 49895;
    i_distance_0054 <= 151784;
    i_distance_0055 <= 235116;
    i_distance_0056 <= 974447;
    i_distance_0057 <= 28796;
    i_distance_0058 <= 333682;
    i_distance_0059 <= 847859;
    i_distance_0060 <= 652274;
    i_distance_0061 <= 1000183;
    i_distance_0062 <= 1004408;
    i_distance_0063 <= 663164;
    correct_answer <= 13410;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 268291;
    i_distance_0001 <= 851079;
    i_distance_0002 <= 898312;
    i_distance_0003 <= 781962;
    i_distance_0004 <= 331661;
    i_distance_0005 <= 993550;
    i_distance_0006 <= 207121;
    i_distance_0007 <= 99986;
    i_distance_0008 <= 99731;
    i_distance_0009 <= 348817;
    i_distance_0010 <= 569365;
    i_distance_0011 <= 342424;
    i_distance_0012 <= 672921;
    i_distance_0013 <= 47002;
    i_distance_0014 <= 653729;
    i_distance_0015 <= 446245;
    i_distance_0016 <= 368551;
    i_distance_0017 <= 977705;
    i_distance_0018 <= 841259;
    i_distance_0019 <= 612652;
    i_distance_0020 <= 445102;
    i_distance_0021 <= 996270;
    i_distance_0022 <= 933808;
    i_distance_0023 <= 192302;
    i_distance_0024 <= 684978;
    i_distance_0025 <= 943026;
    i_distance_0026 <= 331059;
    i_distance_0027 <= 114870;
    i_distance_0028 <= 498999;
    i_distance_0029 <= 653888;
    i_distance_0030 <= 841409;
    i_distance_0031 <= 302784;
    i_distance_0032 <= 1007042;
    i_distance_0033 <= 551492;
    i_distance_0034 <= 413895;
    i_distance_0035 <= 843721;
    i_distance_0036 <= 634573;
    i_distance_0037 <= 219854;
    i_distance_0038 <= 355535;
    i_distance_0039 <= 570703;
    i_distance_0040 <= 68176;
    i_distance_0041 <= 1010902;
    i_distance_0042 <= 436951;
    i_distance_0043 <= 273623;
    i_distance_0044 <= 242905;
    i_distance_0045 <= 956379;
    i_distance_0046 <= 693980;
    i_distance_0047 <= 861;
    i_distance_0048 <= 141532;
    i_distance_0049 <= 255455;
    i_distance_0050 <= 686430;
    i_distance_0051 <= 825953;
    i_distance_0052 <= 863458;
    i_distance_0053 <= 740606;
    i_distance_0054 <= 531175;
    i_distance_0055 <= 482412;
    i_distance_0056 <= 124781;
    i_distance_0057 <= 934256;
    i_distance_0058 <= 182257;
    i_distance_0059 <= 717298;
    i_distance_0060 <= 242802;
    i_distance_0061 <= 651764;
    i_distance_0062 <= 608374;
    i_distance_0063 <= 987390;
    correct_answer <= 861;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 22145;
    i_distance_0001 <= 179971;
    i_distance_0002 <= 722308;
    i_distance_0003 <= 795397;
    i_distance_0004 <= 987398;
    i_distance_0005 <= 663307;
    i_distance_0006 <= 962446;
    i_distance_0007 <= 899857;
    i_distance_0008 <= 731281;
    i_distance_0009 <= 556948;
    i_distance_0010 <= 295963;
    i_distance_0011 <= 823196;
    i_distance_0012 <= 536098;
    i_distance_0013 <= 509347;
    i_distance_0014 <= 974887;
    i_distance_0015 <= 883501;
    i_distance_0016 <= 641966;
    i_distance_0017 <= 866863;
    i_distance_0018 <= 366384;
    i_distance_0019 <= 806321;
    i_distance_0020 <= 215347;
    i_distance_0021 <= 756403;
    i_distance_0022 <= 731445;
    i_distance_0023 <= 981557;
    i_distance_0024 <= 298165;
    i_distance_0025 <= 672057;
    i_distance_0026 <= 718269;
    i_distance_0027 <= 172222;
    i_distance_0028 <= 641599;
    i_distance_0029 <= 1984;
    i_distance_0030 <= 581313;
    i_distance_0031 <= 197183;
    i_distance_0032 <= 806593;
    i_distance_0033 <= 368708;
    i_distance_0034 <= 548037;
    i_distance_0035 <= 942910;
    i_distance_0036 <= 951625;
    i_distance_0037 <= 106570;
    i_distance_0038 <= 945101;
    i_distance_0039 <= 366288;
    i_distance_0040 <= 1009873;
    i_distance_0041 <= 921170;
    i_distance_0042 <= 43859;
    i_distance_0043 <= 400340;
    i_distance_0044 <= 36433;
    i_distance_0045 <= 735321;
    i_distance_0046 <= 705241;
    i_distance_0047 <= 1001178;
    i_distance_0048 <= 116570;
    i_distance_0049 <= 651869;
    i_distance_0050 <= 345052;
    i_distance_0051 <= 551641;
    i_distance_0052 <= 429668;
    i_distance_0053 <= 936293;
    i_distance_0054 <= 619238;
    i_distance_0055 <= 165095;
    i_distance_0056 <= 412010;
    i_distance_0057 <= 865904;
    i_distance_0058 <= 636401;
    i_distance_0059 <= 526450;
    i_distance_0060 <= 294132;
    i_distance_0061 <= 662133;
    i_distance_0062 <= 277495;
    i_distance_0063 <= 626940;
    correct_answer <= 1984;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 854018;
    i_distance_0001 <= 396292;
    i_distance_0002 <= 444292;
    i_distance_0003 <= 264072;
    i_distance_0004 <= 206217;
    i_distance_0005 <= 583433;
    i_distance_0006 <= 151178;
    i_distance_0007 <= 1037580;
    i_distance_0008 <= 312845;
    i_distance_0009 <= 762254;
    i_distance_0010 <= 886030;
    i_distance_0011 <= 816012;
    i_distance_0012 <= 490003;
    i_distance_0013 <= 813715;
    i_distance_0014 <= 900499;
    i_distance_0015 <= 146579;
    i_distance_0016 <= 997780;
    i_distance_0017 <= 711191;
    i_distance_0018 <= 267289;
    i_distance_0019 <= 219543;
    i_distance_0020 <= 209047;
    i_distance_0021 <= 390300;
    i_distance_0022 <= 561693;
    i_distance_0023 <= 417439;
    i_distance_0024 <= 371105;
    i_distance_0025 <= 109729;
    i_distance_0026 <= 457251;
    i_distance_0027 <= 578596;
    i_distance_0028 <= 1007269;
    i_distance_0029 <= 184614;
    i_distance_0030 <= 340265;
    i_distance_0031 <= 958634;
    i_distance_0032 <= 819243;
    i_distance_0033 <= 832306;
    i_distance_0034 <= 320692;
    i_distance_0035 <= 556341;
    i_distance_0036 <= 574646;
    i_distance_0037 <= 622134;
    i_distance_0038 <= 404666;
    i_distance_0039 <= 934204;
    i_distance_0040 <= 704326;
    i_distance_0041 <= 446155;
    i_distance_0042 <= 352209;
    i_distance_0043 <= 534738;
    i_distance_0044 <= 80721;
    i_distance_0045 <= 1025236;
    i_distance_0046 <= 368214;
    i_distance_0047 <= 766427;
    i_distance_0048 <= 560349;
    i_distance_0049 <= 247646;
    i_distance_0050 <= 330846;
    i_distance_0051 <= 36575;
    i_distance_0052 <= 834526;
    i_distance_0053 <= 216542;
    i_distance_0054 <= 579043;
    i_distance_0055 <= 1027303;
    i_distance_0056 <= 345330;
    i_distance_0057 <= 229622;
    i_distance_0058 <= 1046136;
    i_distance_0059 <= 559225;
    i_distance_0060 <= 384250;
    i_distance_0061 <= 844541;
    i_distance_0062 <= 953470;
    i_distance_0063 <= 615935;
    correct_answer <= 36575;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 874625;
    i_distance_0001 <= 993925;
    i_distance_0002 <= 537350;
    i_distance_0003 <= 128265;
    i_distance_0004 <= 671371;
    i_distance_0005 <= 80268;
    i_distance_0006 <= 735375;
    i_distance_0007 <= 529300;
    i_distance_0008 <= 791702;
    i_distance_0009 <= 180760;
    i_distance_0010 <= 209692;
    i_distance_0011 <= 549020;
    i_distance_0012 <= 951967;
    i_distance_0013 <= 557727;
    i_distance_0014 <= 418850;
    i_distance_0015 <= 443049;
    i_distance_0016 <= 758442;
    i_distance_0017 <= 324780;
    i_distance_0018 <= 642350;
    i_distance_0019 <= 89007;
    i_distance_0020 <= 988592;
    i_distance_0021 <= 142256;
    i_distance_0022 <= 731387;
    i_distance_0023 <= 751667;
    i_distance_0024 <= 883123;
    i_distance_0025 <= 898611;
    i_distance_0026 <= 697398;
    i_distance_0027 <= 757687;
    i_distance_0028 <= 782136;
    i_distance_0029 <= 252855;
    i_distance_0030 <= 919226;
    i_distance_0031 <= 671036;
    i_distance_0032 <= 556989;
    i_distance_0033 <= 974656;
    i_distance_0034 <= 929217;
    i_distance_0035 <= 114256;
    i_distance_0036 <= 3538;
    i_distance_0037 <= 402775;
    i_distance_0038 <= 945624;
    i_distance_0039 <= 40920;
    i_distance_0040 <= 774745;
    i_distance_0041 <= 937176;
    i_distance_0042 <= 86874;
    i_distance_0043 <= 804959;
    i_distance_0044 <= 777183;
    i_distance_0045 <= 290657;
    i_distance_0046 <= 32095;
    i_distance_0047 <= 97663;
    i_distance_0048 <= 335849;
    i_distance_0049 <= 554601;
    i_distance_0050 <= 245740;
    i_distance_0051 <= 712556;
    i_distance_0052 <= 553839;
    i_distance_0053 <= 906992;
    i_distance_0054 <= 1777;
    i_distance_0055 <= 680946;
    i_distance_0056 <= 466161;
    i_distance_0057 <= 982389;
    i_distance_0058 <= 522486;
    i_distance_0059 <= 515447;
    i_distance_0060 <= 838777;
    i_distance_0061 <= 741243;
    i_distance_0062 <= 604030;
    i_distance_0063 <= 803839;
    correct_answer <= 1777;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 112130;
    i_distance_0001 <= 1017730;
    i_distance_0002 <= 223238;
    i_distance_0003 <= 732300;
    i_distance_0004 <= 970005;
    i_distance_0005 <= 312214;
    i_distance_0006 <= 95769;
    i_distance_0007 <= 326809;
    i_distance_0008 <= 379545;
    i_distance_0009 <= 303132;
    i_distance_0010 <= 536733;
    i_distance_0011 <= 1032089;
    i_distance_0012 <= 657951;
    i_distance_0013 <= 1024160;
    i_distance_0014 <= 174628;
    i_distance_0015 <= 845349;
    i_distance_0016 <= 832933;
    i_distance_0017 <= 645286;
    i_distance_0018 <= 923688;
    i_distance_0019 <= 617512;
    i_distance_0020 <= 633003;
    i_distance_0021 <= 659116;
    i_distance_0022 <= 47917;
    i_distance_0023 <= 737707;
    i_distance_0024 <= 373165;
    i_distance_0025 <= 529196;
    i_distance_0026 <= 560050;
    i_distance_0027 <= 116284;
    i_distance_0028 <= 832061;
    i_distance_0029 <= 935998;
    i_distance_0030 <= 1007935;
    i_distance_0031 <= 856384;
    i_distance_0032 <= 82241;
    i_distance_0033 <= 713154;
    i_distance_0034 <= 299971;
    i_distance_0035 <= 929345;
    i_distance_0036 <= 502348;
    i_distance_0037 <= 417871;
    i_distance_0038 <= 684752;
    i_distance_0039 <= 695248;
    i_distance_0040 <= 1041744;
    i_distance_0041 <= 149587;
    i_distance_0042 <= 58581;
    i_distance_0043 <= 569047;
    i_distance_0044 <= 164696;
    i_distance_0045 <= 395355;
    i_distance_0046 <= 198621;
    i_distance_0047 <= 30817;
    i_distance_0048 <= 1012451;
    i_distance_0049 <= 437093;
    i_distance_0050 <= 455398;
    i_distance_0051 <= 85991;
    i_distance_0052 <= 511722;
    i_distance_0053 <= 40428;
    i_distance_0054 <= 328430;
    i_distance_0055 <= 248302;
    i_distance_0056 <= 262896;
    i_distance_0057 <= 864243;
    i_distance_0058 <= 967027;
    i_distance_0059 <= 11251;
    i_distance_0060 <= 391412;
    i_distance_0061 <= 81655;
    i_distance_0062 <= 901497;
    i_distance_0063 <= 36860;
    correct_answer <= 11251;
    sync_wait_rising(clk, 10);

    i_distance_0000 <= 72834;
    i_distance_0001 <= 650500;
    i_distance_0002 <= 174084;
    i_distance_0003 <= 169349;
    i_distance_0004 <= 146696;
    i_distance_0005 <= 287884;
    i_distance_0006 <= 747407;
    i_distance_0007 <= 480655;
    i_distance_0008 <= 890129;
    i_distance_0009 <= 215443;
    i_distance_0010 <= 81177;
    i_distance_0011 <= 5529;
    i_distance_0012 <= 282010;
    i_distance_0013 <= 569626;
    i_distance_0014 <= 718626;
    i_distance_0015 <= 278053;
    i_distance_0016 <= 383783;
    i_distance_0017 <= 530219;
    i_distance_0018 <= 281516;
    i_distance_0019 <= 841773;
    i_distance_0020 <= 874544;
    i_distance_0021 <= 693680;
    i_distance_0022 <= 578225;
    i_distance_0023 <= 305587;
    i_distance_0024 <= 119091;
    i_distance_0025 <= 866742;
    i_distance_0026 <= 773050;
    i_distance_0027 <= 602811;
    i_distance_0028 <= 304445;
    i_distance_0029 <= 720189;
    i_distance_0030 <= 291904;
    i_distance_0031 <= 898753;
    i_distance_0032 <= 470466;
    i_distance_0033 <= 9923;
    i_distance_0034 <= 57157;
    i_distance_0035 <= 608838;
    i_distance_0036 <= 297032;
    i_distance_0037 <= 455627;
    i_distance_0038 <= 42956;
    i_distance_0039 <= 520267;
    i_distance_0040 <= 496079;
    i_distance_0041 <= 978512;
    i_distance_0042 <= 22737;
    i_distance_0043 <= 543825;
    i_distance_0044 <= 778191;
    i_distance_0045 <= 193620;
    i_distance_0046 <= 590810;
    i_distance_0047 <= 400348;
    i_distance_0048 <= 863837;
    i_distance_0049 <= 546145;
    i_distance_0050 <= 985058;
    i_distance_0051 <= 815457;
    i_distance_0052 <= 466148;
    i_distance_0053 <= 154081;
    i_distance_0054 <= 638567;
    i_distance_0055 <= 57193;
    i_distance_0056 <= 524778;
    i_distance_0057 <= 26218;
    i_distance_0058 <= 691310;
    i_distance_0059 <= 269552;
    i_distance_0060 <= 747637;
    i_distance_0061 <= 440695;
    i_distance_0062 <= 281340;
    i_distance_0063 <= 816894;
    correct_answer <= 5529;
    sync_wait_rising(clk, 10);
    
    sync_wait_rising(clk, 100);
    sim_done <= '1';
    wait;
end process;




----------------------------------------------------------------------------------------------------
--                                        Unit Under Test
----------------------------------------------------------------------------------------------------
UUT: MinFunction_0064 port map (
    clk => clk,
    rst => rst,
    i_soft_rst => i_soft_rst,
    i_distance_0000 => i_distance_0000,
    i_distance_0001 => i_distance_0001,
    i_distance_0002 => i_distance_0002,
    i_distance_0003 => i_distance_0003,
    i_distance_0004 => i_distance_0004,
    i_distance_0005 => i_distance_0005,
    i_distance_0006 => i_distance_0006,
    i_distance_0007 => i_distance_0007,
    i_distance_0008 => i_distance_0008,
    i_distance_0009 => i_distance_0009,
    i_distance_0010 => i_distance_0010,
    i_distance_0011 => i_distance_0011,
    i_distance_0012 => i_distance_0012,
    i_distance_0013 => i_distance_0013,
    i_distance_0014 => i_distance_0014,
    i_distance_0015 => i_distance_0015,
    i_distance_0016 => i_distance_0016,
    i_distance_0017 => i_distance_0017,
    i_distance_0018 => i_distance_0018,
    i_distance_0019 => i_distance_0019,
    i_distance_0020 => i_distance_0020,
    i_distance_0021 => i_distance_0021,
    i_distance_0022 => i_distance_0022,
    i_distance_0023 => i_distance_0023,
    i_distance_0024 => i_distance_0024,
    i_distance_0025 => i_distance_0025,
    i_distance_0026 => i_distance_0026,
    i_distance_0027 => i_distance_0027,
    i_distance_0028 => i_distance_0028,
    i_distance_0029 => i_distance_0029,
    i_distance_0030 => i_distance_0030,
    i_distance_0031 => i_distance_0031,
    i_distance_0032 => i_distance_0032,
    i_distance_0033 => i_distance_0033,
    i_distance_0034 => i_distance_0034,
    i_distance_0035 => i_distance_0035,
    i_distance_0036 => i_distance_0036,
    i_distance_0037 => i_distance_0037,
    i_distance_0038 => i_distance_0038,
    i_distance_0039 => i_distance_0039,
    i_distance_0040 => i_distance_0040,
    i_distance_0041 => i_distance_0041,
    i_distance_0042 => i_distance_0042,
    i_distance_0043 => i_distance_0043,
    i_distance_0044 => i_distance_0044,
    i_distance_0045 => i_distance_0045,
    i_distance_0046 => i_distance_0046,
    i_distance_0047 => i_distance_0047,
    i_distance_0048 => i_distance_0048,
    i_distance_0049 => i_distance_0049,
    i_distance_0050 => i_distance_0050,
    i_distance_0051 => i_distance_0051,
    i_distance_0052 => i_distance_0052,
    i_distance_0053 => i_distance_0053,
    i_distance_0054 => i_distance_0054,
    i_distance_0055 => i_distance_0055,
    i_distance_0056 => i_distance_0056,
    i_distance_0057 => i_distance_0057,
    i_distance_0058 => i_distance_0058,
    i_distance_0059 => i_distance_0059,
    i_distance_0060 => i_distance_0060,
    i_distance_0061 => i_distance_0061,
    i_distance_0062 => i_distance_0062,
    i_distance_0063 => i_distance_0063,
    o_min => o_min,
    o_latency => o_latency
);


end architecture behavioral_MinFunction_0064_tb;


