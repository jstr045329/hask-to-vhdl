library ieee;
use ieee.std_logic_1164.all;


entity count1s is
    generic (
        use_async_reset : std_logic := '1'
    );
    port (
        clk : in std_logic;
        reset : in std_logic;
        a0 : in std_logic := '0';
        a1 : in std_logic := '0';
        a2 : in std_logic := '0';
        a3 : in std_logic := '0';
        a4 : in std_logic := '0';
        a5 : in std_logic := '0';
        a6 : in std_logic := '0';
        a7 : in std_logic := '0';
        q : out std_logic_vector(3 downto 0)
    );
end count1s;


architecture behavioral_count1s of count1s is

signal agg : std_logic_vector(3 downto 0);

function count_bits(
    x : std_logic_vector(7 downto 0)
    ) return std_logic_vector is
variable y : std_logic_vector(3 downto 0);
begin
    y := (others => '0');
    case x is
    when "00000000" =>
        y := "0000";
    when "00000001" =>
        y := "0001";
    when "00000010" =>
        y := "0001";
    when "00000011" =>
        y := "0010";
    when "00000100" =>
        y := "0001";
    when "00000101" =>
        y := "0010";
    when "00000110" =>
        y := "0010";
    when "00000111" =>
        y := "0011";
    when "00001000" =>
        y := "0001";
    when "00001001" =>
        y := "0010";
    when "00001010" =>
        y := "0010";
    when "00001011" =>
        y := "0011";
    when "00001100" =>
        y := "0010";
    when "00001101" =>
        y := "0011";
    when "00001110" =>
        y := "0011";
    when "00001111" =>
        y := "0100";
    when "00010000" =>
        y := "0001";
    when "00010001" =>
        y := "0010";
    when "00010010" =>
        y := "0010";
    when "00010011" =>
        y := "0011";
    when "00010100" =>
        y := "0010";
    when "00010101" =>
        y := "0011";
    when "00010110" =>
        y := "0011";
    when "00010111" =>
        y := "0100";
    when "00011000" =>
        y := "0010";
    when "00011001" =>
        y := "0011";
    when "00011010" =>
        y := "0011";
    when "00011011" =>
        y := "0100";
    when "00011100" =>
        y := "0011";
    when "00011101" =>
        y := "0100";
    when "00011110" =>
        y := "0100";
    when "00011111" =>
        y := "0101";
    when "00100000" =>
        y := "0001";
    when "00100001" =>
        y := "0010";
    when "00100010" =>
        y := "0010";
    when "00100011" =>
        y := "0011";
    when "00100100" =>
        y := "0010";
    when "00100101" =>
        y := "0011";
    when "00100110" =>
        y := "0011";
    when "00100111" =>
        y := "0100";
    when "00101000" =>
        y := "0010";
    when "00101001" =>
        y := "0011";
    when "00101010" =>
        y := "0011";
    when "00101011" =>
        y := "0100";
    when "00101100" =>
        y := "0011";
    when "00101101" =>
        y := "0100";
    when "00101110" =>
        y := "0100";
    when "00101111" =>
        y := "0101";
    when "00110000" =>
        y := "0010";
    when "00110001" =>
        y := "0011";
    when "00110010" =>
        y := "0011";
    when "00110011" =>
        y := "0100";
    when "00110100" =>
        y := "0011";
    when "00110101" =>
        y := "0100";
    when "00110110" =>
        y := "0100";
    when "00110111" =>
        y := "0101";
    when "00111000" =>
        y := "0011";
    when "00111001" =>
        y := "0100";
    when "00111010" =>
        y := "0100";
    when "00111011" =>
        y := "0101";
    when "00111100" =>
        y := "0100";
    when "00111101" =>
        y := "0101";
    when "00111110" =>
        y := "0101";
    when "00111111" =>
        y := "0110";
    when "01000000" =>
        y := "0001";
    when "01000001" =>
        y := "0010";
    when "01000010" =>
        y := "0010";
    when "01000011" =>
        y := "0011";
    when "01000100" =>
        y := "0010";
    when "01000101" =>
        y := "0011";
    when "01000110" =>
        y := "0011";
    when "01000111" =>
        y := "0100";
    when "01001000" =>
        y := "0010";
    when "01001001" =>
        y := "0011";
    when "01001010" =>
        y := "0011";
    when "01001011" =>
        y := "0100";
    when "01001100" =>
        y := "0011";
    when "01001101" =>
        y := "0100";
    when "01001110" =>
        y := "0100";
    when "01001111" =>
        y := "0101";
    when "01010000" =>
        y := "0010";
    when "01010001" =>
        y := "0011";
    when "01010010" =>
        y := "0011";
    when "01010011" =>
        y := "0100";
    when "01010100" =>
        y := "0011";
    when "01010101" =>
        y := "0100";
    when "01010110" =>
        y := "0100";
    when "01010111" =>
        y := "0101";
    when "01011000" =>
        y := "0011";
    when "01011001" =>
        y := "0100";
    when "01011010" =>
        y := "0100";
    when "01011011" =>
        y := "0101";
    when "01011100" =>
        y := "0100";
    when "01011101" =>
        y := "0101";
    when "01011110" =>
        y := "0101";
    when "01011111" =>
        y := "0110";
    when "01100000" =>
        y := "0010";
    when "01100001" =>
        y := "0011";
    when "01100010" =>
        y := "0011";
    when "01100011" =>
        y := "0100";
    when "01100100" =>
        y := "0011";
    when "01100101" =>
        y := "0100";
    when "01100110" =>
        y := "0100";
    when "01100111" =>
        y := "0101";
    when "01101000" =>
        y := "0011";
    when "01101001" =>
        y := "0100";
    when "01101010" =>
        y := "0100";
    when "01101011" =>
        y := "0101";
    when "01101100" =>
        y := "0100";
    when "01101101" =>
        y := "0101";
    when "01101110" =>
        y := "0101";
    when "01101111" =>
        y := "0110";
    when "01110000" =>
        y := "0011";
    when "01110001" =>
        y := "0100";
    when "01110010" =>
        y := "0100";
    when "01110011" =>
        y := "0101";
    when "01110100" =>
        y := "0100";
    when "01110101" =>
        y := "0101";
    when "01110110" =>
        y := "0101";
    when "01110111" =>
        y := "0110";
    when "01111000" =>
        y := "0100";
    when "01111001" =>
        y := "0101";
    when "01111010" =>
        y := "0101";
    when "01111011" =>
        y := "0110";
    when "01111100" =>
        y := "0101";
    when "01111101" =>
        y := "0110";
    when "01111110" =>
        y := "0110";
    when "01111111" =>
        y := "0111";
    when "10000000" =>
        y := "0001";
    when "10000001" =>
        y := "0010";
    when "10000010" =>
        y := "0010";
    when "10000011" =>
        y := "0011";
    when "10000100" =>
        y := "0010";
    when "10000101" =>
        y := "0011";
    when "10000110" =>
        y := "0011";
    when "10000111" =>
        y := "0100";
    when "10001000" =>
        y := "0010";
    when "10001001" =>
        y := "0011";
    when "10001010" =>
        y := "0011";
    when "10001011" =>
        y := "0100";
    when "10001100" =>
        y := "0011";
    when "10001101" =>
        y := "0100";
    when "10001110" =>
        y := "0100";
    when "10001111" =>
        y := "0101";
    when "10010000" =>
        y := "0010";
    when "10010001" =>
        y := "0011";
    when "10010010" =>
        y := "0011";
    when "10010011" =>
        y := "0100";
    when "10010100" =>
        y := "0011";
    when "10010101" =>
        y := "0100";
    when "10010110" =>
        y := "0100";
    when "10010111" =>
        y := "0101";
    when "10011000" =>
        y := "0011";
    when "10011001" =>
        y := "0100";
    when "10011010" =>
        y := "0100";
    when "10011011" =>
        y := "0101";
    when "10011100" =>
        y := "0100";
    when "10011101" =>
        y := "0101";
    when "10011110" =>
        y := "0101";
    when "10011111" =>
        y := "0110";
    when "10100000" =>
        y := "0010";
    when "10100001" =>
        y := "0011";
    when "10100010" =>
        y := "0011";
    when "10100011" =>
        y := "0100";
    when "10100100" =>
        y := "0011";
    when "10100101" =>
        y := "0100";
    when "10100110" =>
        y := "0100";
    when "10100111" =>
        y := "0101";
    when "10101000" =>
        y := "0011";
    when "10101001" =>
        y := "0100";
    when "10101010" =>
        y := "0100";
    when "10101011" =>
        y := "0101";
    when "10101100" =>
        y := "0100";
    when "10101101" =>
        y := "0101";
    when "10101110" =>
        y := "0101";
    when "10101111" =>
        y := "0110";
    when "10110000" =>
        y := "0011";
    when "10110001" =>
        y := "0100";
    when "10110010" =>
        y := "0100";
    when "10110011" =>
        y := "0101";
    when "10110100" =>
        y := "0100";
    when "10110101" =>
        y := "0101";
    when "10110110" =>
        y := "0101";
    when "10110111" =>
        y := "0110";
    when "10111000" =>
        y := "0100";
    when "10111001" =>
        y := "0101";
    when "10111010" =>
        y := "0101";
    when "10111011" =>
        y := "0110";
    when "10111100" =>
        y := "0101";
    when "10111101" =>
        y := "0110";
    when "10111110" =>
        y := "0110";
    when "10111111" =>
        y := "0111";
    when "11000000" =>
        y := "0010";
    when "11000001" =>
        y := "0011";
    when "11000010" =>
        y := "0011";
    when "11000011" =>
        y := "0100";
    when "11000100" =>
        y := "0011";
    when "11000101" =>
        y := "0100";
    when "11000110" =>
        y := "0100";
    when "11000111" =>
        y := "0101";
    when "11001000" =>
        y := "0011";
    when "11001001" =>
        y := "0100";
    when "11001010" =>
        y := "0100";
    when "11001011" =>
        y := "0101";
    when "11001100" =>
        y := "0100";
    when "11001101" =>
        y := "0101";
    when "11001110" =>
        y := "0101";
    when "11001111" =>
        y := "0110";
    when "11010000" =>
        y := "0011";
    when "11010001" =>
        y := "0100";
    when "11010010" =>
        y := "0100";
    when "11010011" =>
        y := "0101";
    when "11010100" =>
        y := "0100";
    when "11010101" =>
        y := "0101";
    when "11010110" =>
        y := "0101";
    when "11010111" =>
        y := "0110";
    when "11011000" =>
        y := "0100";
    when "11011001" =>
        y := "0101";
    when "11011010" =>
        y := "0101";
    when "11011011" =>
        y := "0110";
    when "11011100" =>
        y := "0101";
    when "11011101" =>
        y := "0110";
    when "11011110" =>
        y := "0110";
    when "11011111" =>
        y := "0111";
    when "11100000" =>
        y := "0011";
    when "11100001" =>
        y := "0100";
    when "11100010" =>
        y := "0100";
    when "11100011" =>
        y := "0101";
    when "11100100" =>
        y := "0100";
    when "11100101" =>
        y := "0101";
    when "11100110" =>
        y := "0101";
    when "11100111" =>
        y := "0110";
    when "11101000" =>
        y := "0100";
    when "11101001" =>
        y := "0101";
    when "11101010" =>
        y := "0101";
    when "11101011" =>
        y := "0110";
    when "11101100" =>
        y := "0101";
    when "11101101" =>
        y := "0110";
    when "11101110" =>
        y := "0110";
    when "11101111" =>
        y := "0111";
    when "11110000" =>
        y := "0100";
    when "11110001" =>
        y := "0101";
    when "11110010" =>
        y := "0101";
    when "11110011" =>
        y := "0110";
    when "11110100" =>
        y := "0101";
    when "11110101" =>
        y := "0110";
    when "11110110" =>
        y := "0110";
    when "11110111" =>
        y := "0111";
    when "11111000" =>
        y := "0101";
    when "11111001" =>
        y := "0110";
    when "11111010" =>
        y := "0110";
    when "11111011" =>
        y := "0111";
    when "11111100" =>
        y := "0110";
    when "11111101" =>
        y := "0111";
    when "11111110" =>
        y := "0111";
    when "11111111" =>
        y := "1000";
    when others =>
        y := (others => '0');
    end case;
    return y;
end function;


begin

agg <= a0 & a1 & a2 & a3 & a4 & a5 & a6 & a7;

USE_ASYNC_RESET_BLOCK: if use_async_reset = '1' generate 
    process(clk, reset)
    begin
        if reset = '1' then
            q <= (others => '0');
        elsif rising_edge(clk) then
            q <= count_bits(agg);
        end if;
    end process;
end generate;

USE_SYNC_RESET_BLOCK: if use_async_reset = '0' generate
    process(clk)
    begin
        if rising_edge(clk) then
            if reset = '1' then
                q <= (others => '0');
            else
                q <= count_bits(agg);
            end if;
        end if;
    end process;
end generate;

end behavioral_count1s;


