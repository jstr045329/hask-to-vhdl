-- <entities_here>

library IEEE;
use IEEE.std_logic_1164.ALL;
use IEEE.numeric_std.ALL;
use work.PowerSetGears.all;


------------------------------------------------------------------------------------------------------------------------
--                                        At Long Last: The Power Set Package 
------------------------------------------------------------------------------------------------------------------------
package PowerSetPkg is

-- <component_declarations_here>

end package PowerSetPkg;


package body PowerSetPkg is
end package body PowerSetPkg;
