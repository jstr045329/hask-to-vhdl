------------------------------------------------------------------------------------------------------------------------
--                        Test Variadic Logic Functions in SingleCyclePipelinedFunctions.vhd 
--
-- This testbench tests functions in the SingleCyclePipelinedFunctions package. Because the UUT's are functions, 
-- not entities, there is no component instantiation at the bottom like there normally is. Instead, there are only 
-- function calls. 
--
------------------------------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.VhdSimToolsPkg.all;
use work.SingleCyclePipelinedFunctions.all;


entity TestVariadicLogicFunctions_tb is
end TestVariadicLogicFunctions_tb;


architecture behavioral_TestVariadicLogicFunctions_tb of TestVariadicLogicFunctions_tb is

signal clk : std_logic := '1';
signal rst : std_logic := '1';

constant clk_per : time := 10 ns;
signal sim_done : std_logic := '0';
signal test_stage : integer := 0;
signal s_clock_cycle_count : integer := 0;
signal s_x : std_logic_vector(255 downto 0);
signal s_and_chain : std_logic_vector(255 downto 0);
signal y_and : std_logic := '0';
signal y_or : std_logic := '0';
signal y_nand : std_logic := '0';
signal y_nor : std_logic := '0';
signal y_xor : std_logic := '0';
signal x_feed : std_logic;

begin


----------------------------------------------------------------------------------------------------
--                                          Boiler Plate
----------------------------------------------------------------------------------------------------
CLOCK_PROCESS: process
begin
    if sim_done = '1' then
        wait;
    else
        wait for clk_per/2;
        clk <= not clk;
    end if;
end process;


----------------------------------------------------------------------------------------------------
--                                       Count Clock Cycles
----------------------------------------------------------------------------------------------------
CLOCK_CYCLE_COUNTER: process(clk)
begin
    if rising_edge(clk) then 
        s_clock_cycle_count <= s_clock_cycle_count + 1;
    end if;
end process;


------------------------------------------------------------------------------------------------------------------------
--                            Stim Process 1: Form The Input Signals Into A Long Pipeline 
------------------------------------------------------------------------------------------------------------------------
STIM_PROCESS_1:process(clk)
begin
    if rising_edge(clk) then 
        if rst = '1' then 
            s_x <= (others => '0');
            s_and_chain <= (others => '1');
        else
            s_x <= x_feed & s_x(255 downto 1);
            s_and_chain <= (not x_feed) & s_and_chain(255 downto 1);
        end if;
    end if;
end process;



------------------------------------------------------------------------------------------------------------------------
--                                   Stim Process 2: Do Normal Stim Process Stuff 
------------------------------------------------------------------------------------------------------------------------
STIM_PROCESS_2: process
begin
    x_feed <= '0';
    test_stage <= 0;
    sync_wait_rising(clk, 10);
    rst <= not rst;
    sync_wait_rising(clk, 10);
    
    -- Strobe the signal that feeds a pulse into the delay line:
    strobe_rising(clk, x_feed);

    -- Let UUT do its thing:
    for i in 0 to 255 loop
        sync_wait_rising(clk, 1);
    end loop;

    -- Test ends here:
    test_stage <= test_stage + 1;
    sync_wait_rising(clk, 100);
    sim_done <= '1';
    wait;
end process;


------------------------------------------------------------------------------------------------------------------------
--                                               Unit Under Test (UUT) 
------------------------------------------------------------------------------------------------------------------------
y_and <= large_and(
    s_and_chain(1),
    s_and_chain(3),
    s_and_chain(5),
    s_and_chain(7),
    s_and_chain(9),
    s_and_chain(11),
    s_and_chain(13),
    s_and_chain(15),
    s_and_chain(17),
    s_and_chain(19),
    s_and_chain(21),
    s_and_chain(23),
    s_and_chain(25),
    s_and_chain(27),
    s_and_chain(29),
    s_and_chain(31),
    s_and_chain(33),
    s_and_chain(35),
    s_and_chain(37),
    s_and_chain(39),
    s_and_chain(41),
    s_and_chain(43),
    s_and_chain(45),
    s_and_chain(47),
    s_and_chain(49),
    s_and_chain(51),
    s_and_chain(53),
    s_and_chain(55),
    s_and_chain(57),
    s_and_chain(59),
    s_and_chain(61),
    s_and_chain(63),
    s_and_chain(65),
    s_and_chain(67),
    s_and_chain(69),
    s_and_chain(71),
    s_and_chain(73),
    s_and_chain(75),
    s_and_chain(77),
    s_and_chain(79),
    s_and_chain(81),
    s_and_chain(83),
    s_and_chain(85),
    s_and_chain(87),
    s_and_chain(89),
    s_and_chain(91),
    s_and_chain(93),
    s_and_chain(95),
    s_and_chain(97),
    s_and_chain(99),
    s_and_chain(101),
    s_and_chain(103),
    s_and_chain(105),
    s_and_chain(107),
    s_and_chain(109),
    s_and_chain(111),
    s_and_chain(113),
    s_and_chain(115),
    s_and_chain(117),
    s_and_chain(119),
    s_and_chain(121),
    s_and_chain(123),
    s_and_chain(125),
    s_and_chain(127),
    s_and_chain(129),
    s_and_chain(131),
    s_and_chain(133),
    s_and_chain(135),
    s_and_chain(137),
    s_and_chain(139),
    s_and_chain(141),
    s_and_chain(143),
    s_and_chain(145),
    s_and_chain(147),
    s_and_chain(149),
    s_and_chain(151),
    s_and_chain(153),
    s_and_chain(155),
    s_and_chain(157),
    s_and_chain(159),
    s_and_chain(161),
    s_and_chain(163),
    s_and_chain(165),
    s_and_chain(167),
    s_and_chain(169),
    s_and_chain(171),
    s_and_chain(173),
    s_and_chain(175),
    s_and_chain(177),
    s_and_chain(179),
    s_and_chain(181),
    s_and_chain(183),
    s_and_chain(185),
    s_and_chain(187),
    s_and_chain(189),
    s_and_chain(191),
    s_and_chain(193),
    s_and_chain(195),
    s_and_chain(197),
    s_and_chain(199),
    s_and_chain(201),
    s_and_chain(203),
    s_and_chain(205),
    s_and_chain(207),
    s_and_chain(209),
    s_and_chain(211),
    s_and_chain(213),
    s_and_chain(215),
    s_and_chain(217),
    s_and_chain(219),
    s_and_chain(221),
    s_and_chain(223),
    s_and_chain(225),
    s_and_chain(227),
    s_and_chain(229),
    s_and_chain(231),
    s_and_chain(233),
    s_and_chain(235),
    s_and_chain(237),
    s_and_chain(239),
    s_and_chain(241),
    s_and_chain(243),
    s_and_chain(245),
    s_and_chain(247),
    s_and_chain(249),
    s_and_chain(251),
    s_and_chain(253),
    s_and_chain(255)
    );



y_or <= large_or(
    s_x(1),
    s_x(3),
    s_x(5),
    s_x(7),
    s_x(9),
    s_x(11),
    s_x(13),
    s_x(15),
    s_x(17),
    s_x(19),
    s_x(21),
    s_x(23),
    s_x(25),
    s_x(27),
    s_x(29),
    s_x(31),
    s_x(33),
    s_x(35),
    s_x(37),
    s_x(39),
    s_x(41),
    s_x(43),
    s_x(45),
    s_x(47),
    s_x(49),
    s_x(51),
    s_x(53),
    s_x(55),
    s_x(57),
    s_x(59),
    s_x(61),
    s_x(63),
    s_x(65),
    s_x(67),
    s_x(69),
    s_x(71),
    s_x(73),
    s_x(75),
    s_x(77),
    s_x(79),
    s_x(81),
    s_x(83),
    s_x(85),
    s_x(87),
    s_x(89),
    s_x(91),
    s_x(93),
    s_x(95),
    s_x(97),
    s_x(99),
    s_x(101),
    s_x(103),
    s_x(105),
    s_x(107),
    s_x(109),
    s_x(111),
    s_x(113),
    s_x(115),
    s_x(117),
    s_x(119),
    s_x(121),
    s_x(123),
    s_x(125),
    s_x(127),
    s_x(129),
    s_x(131),
    s_x(133),
    s_x(135),
    s_x(137),
    s_x(139),
    s_x(141),
    s_x(143),
    s_x(145),
    s_x(147),
    s_x(149),
    s_x(151),
    s_x(153),
    s_x(155),
    s_x(157),
    s_x(159),
    s_x(161),
    s_x(163),
    s_x(165),
    s_x(167),
    s_x(169),
    s_x(171),
    s_x(173),
    s_x(175),
    s_x(177),
    s_x(179),
    s_x(181),
    s_x(183),
    s_x(185),
    s_x(187),
    s_x(189),
    s_x(191),
    s_x(193),
    s_x(195),
    s_x(197),
    s_x(199),
    s_x(201),
    s_x(203),
    s_x(205),
    s_x(207),
    s_x(209),
    s_x(211),
    s_x(213),
    s_x(215),
    s_x(217),
    s_x(219),
    s_x(221),
    s_x(223),
    s_x(225),
    s_x(227),
    s_x(229),
    s_x(231),
    s_x(233),
    s_x(235),
    s_x(237),
    s_x(239),
    s_x(241),
    s_x(243),
    s_x(245),
    s_x(247),
    s_x(249),
    s_x(251),
    s_x(253),
    s_x(255)
    );


y_nand <= large_nand(
    s_and_chain(1),
    s_and_chain(3),
    s_and_chain(5),
    s_and_chain(7),
    s_and_chain(9),
    s_and_chain(11),
    s_and_chain(13),
    s_and_chain(15),
    s_and_chain(17),
    s_and_chain(19),
    s_and_chain(21),
    s_and_chain(23),
    s_and_chain(25),
    s_and_chain(27),
    s_and_chain(29),
    s_and_chain(31),
    s_and_chain(33),
    s_and_chain(35),
    s_and_chain(37),
    s_and_chain(39),
    s_and_chain(41),
    s_and_chain(43),
    s_and_chain(45),
    s_and_chain(47),
    s_and_chain(49),
    s_and_chain(51),
    s_and_chain(53),
    s_and_chain(55),
    s_and_chain(57),
    s_and_chain(59),
    s_and_chain(61),
    s_and_chain(63),
    s_and_chain(65),
    s_and_chain(67),
    s_and_chain(69),
    s_and_chain(71),
    s_and_chain(73),
    s_and_chain(75),
    s_and_chain(77),
    s_and_chain(79),
    s_and_chain(81),
    s_and_chain(83),
    s_and_chain(85),
    s_and_chain(87),
    s_and_chain(89),
    s_and_chain(91),
    s_and_chain(93),
    s_and_chain(95),
    s_and_chain(97),
    s_and_chain(99),
    s_and_chain(101),
    s_and_chain(103),
    s_and_chain(105),
    s_and_chain(107),
    s_and_chain(109),
    s_and_chain(111),
    s_and_chain(113),
    s_and_chain(115),
    s_and_chain(117),
    s_and_chain(119),
    s_and_chain(121),
    s_and_chain(123),
    s_and_chain(125),
    s_and_chain(127),
    s_and_chain(129),
    s_and_chain(131),
    s_and_chain(133),
    s_and_chain(135),
    s_and_chain(137),
    s_and_chain(139),
    s_and_chain(141),
    s_and_chain(143),
    s_and_chain(145),
    s_and_chain(147),
    s_and_chain(149),
    s_and_chain(151),
    s_and_chain(153),
    s_and_chain(155),
    s_and_chain(157),
    s_and_chain(159),
    s_and_chain(161),
    s_and_chain(163),
    s_and_chain(165),
    s_and_chain(167),
    s_and_chain(169),
    s_and_chain(171),
    s_and_chain(173),
    s_and_chain(175),
    s_and_chain(177),
    s_and_chain(179),
    s_and_chain(181),
    s_and_chain(183),
    s_and_chain(185),
    s_and_chain(187),
    s_and_chain(189),
    s_and_chain(191),
    s_and_chain(193),
    s_and_chain(195),
    s_and_chain(197),
    s_and_chain(199),
    s_and_chain(201),
    s_and_chain(203),
    s_and_chain(205),
    s_and_chain(207),
    s_and_chain(209),
    s_and_chain(211),
    s_and_chain(213),
    s_and_chain(215),
    s_and_chain(217),
    s_and_chain(219),
    s_and_chain(221),
    s_and_chain(223),
    s_and_chain(225),
    s_and_chain(227),
    s_and_chain(229),
    s_and_chain(231),
    s_and_chain(233),
    s_and_chain(235),
    s_and_chain(237),
    s_and_chain(239),
    s_and_chain(241),
    s_and_chain(243),
    s_and_chain(245),
    s_and_chain(247),
    s_and_chain(249),
    s_and_chain(251),
    s_and_chain(253),
    s_and_chain(255)
    );


y_nor <= large_nor(
    s_x(1),
    s_x(3),
    s_x(5),
    s_x(7),
    s_x(9),
    s_x(11),
    s_x(13),
    s_x(15),
    s_x(17),
    s_x(19),
    s_x(21),
    s_x(23),
    s_x(25),
    s_x(27),
    s_x(29),
    s_x(31),
    s_x(33),
    s_x(35),
    s_x(37),
    s_x(39),
    s_x(41),
    s_x(43),
    s_x(45),
    s_x(47),
    s_x(49),
    s_x(51),
    s_x(53),
    s_x(55),
    s_x(57),
    s_x(59),
    s_x(61),
    s_x(63),
    s_x(65),
    s_x(67),
    s_x(69),
    s_x(71),
    s_x(73),
    s_x(75),
    s_x(77),
    s_x(79),
    s_x(81),
    s_x(83),
    s_x(85),
    s_x(87),
    s_x(89),
    s_x(91),
    s_x(93),
    s_x(95),
    s_x(97),
    s_x(99),
    s_x(101),
    s_x(103),
    s_x(105),
    s_x(107),
    s_x(109),
    s_x(111),
    s_x(113),
    s_x(115),
    s_x(117),
    s_x(119),
    s_x(121),
    s_x(123),
    s_x(125),
    s_x(127),
    s_x(129),
    s_x(131),
    s_x(133),
    s_x(135),
    s_x(137),
    s_x(139),
    s_x(141),
    s_x(143),
    s_x(145),
    s_x(147),
    s_x(149),
    s_x(151),
    s_x(153),
    s_x(155),
    s_x(157),
    s_x(159),
    s_x(161),
    s_x(163),
    s_x(165),
    s_x(167),
    s_x(169),
    s_x(171),
    s_x(173),
    s_x(175),
    s_x(177),
    s_x(179),
    s_x(181),
    s_x(183),
    s_x(185),
    s_x(187),
    s_x(189),
    s_x(191),
    s_x(193),
    s_x(195),
    s_x(197),
    s_x(199),
    s_x(201),
    s_x(203),
    s_x(205),
    s_x(207),
    s_x(209),
    s_x(211),
    s_x(213),
    s_x(215),
    s_x(217),
    s_x(219),
    s_x(221),
    s_x(223),
    s_x(225),
    s_x(227),
    s_x(229),
    s_x(231),
    s_x(233),
    s_x(235),
    s_x(237),
    s_x(239),
    s_x(241),
    s_x(243),
    s_x(245),
    s_x(247),
    s_x(249),
    s_x(251),
    s_x(253),
    s_x(255)
    );


y_xor <= large_xor(
    s_x(1),
    s_x(3),
    s_x(5),
    s_x(7),
    s_x(9),
    s_x(11),
    s_x(13),
    s_x(15),
    s_x(17),
    s_x(19),
    s_x(21),
    s_x(23),
    s_x(25),
    s_x(27),
    s_x(29),
    s_x(31),
    s_x(33),
    s_x(35),
    s_x(37),
    s_x(39),
    s_x(41),
    s_x(43),
    s_x(45),
    s_x(47),
    s_x(49),
    s_x(51),
    s_x(53),
    s_x(55),
    s_x(57),
    s_x(59),
    s_x(61),
    s_x(63),
    s_x(65),
    s_x(67),
    s_x(69),
    s_x(71),
    s_x(73),
    s_x(75),
    s_x(77),
    s_x(79),
    s_x(81),
    s_x(83),
    s_x(85),
    s_x(87),
    s_x(89),
    s_x(91),
    s_x(93),
    s_x(95),
    s_x(97),
    s_x(99),
    s_x(101),
    s_x(103),
    s_x(105),
    s_x(107),
    s_x(109),
    s_x(111),
    s_x(113),
    s_x(115),
    s_x(117),
    s_x(119),
    s_x(121),
    s_x(123),
    s_x(125),
    s_x(127),
    s_x(129),
    s_x(131),
    s_x(133),
    s_x(135),
    s_x(137),
    s_x(139),
    s_x(141),
    s_x(143),
    s_x(145),
    s_x(147),
    s_x(149),
    s_x(151),
    s_x(153),
    s_x(155),
    s_x(157),
    s_x(159),
    s_x(161),
    s_x(163),
    s_x(165),
    s_x(167),
    s_x(169),
    s_x(171),
    s_x(173),
    s_x(175),
    s_x(177),
    s_x(179),
    s_x(181),
    s_x(183),
    s_x(185),
    s_x(187),
    s_x(189),
    s_x(191),
    s_x(193),
    s_x(195),
    s_x(197),
    s_x(199),
    s_x(201),
    s_x(203),
    s_x(205),
    s_x(207),
    s_x(209),
    s_x(211),
    s_x(213),
    s_x(215),
    s_x(217),
    s_x(219),
    s_x(221),
    s_x(223),
    s_x(225),
    s_x(227),
    s_x(229),
    s_x(231),
    s_x(233),
    s_x(235),
    s_x(237),
    s_x(239),
    s_x(241),
    s_x(243),
    s_x(245),
    s_x(247),
    s_x(249),
    s_x(251),
    s_x(253),
    s_x(255)
    );


end architecture behavioral_TestVariadicLogicFunctions_tb;


