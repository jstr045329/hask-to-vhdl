library IEEE;
use IEEE.std_logic_1164.ALL;
use IEEE.numeric_std.ALL;
use work.RegisteredGatesPkg.all;


entity ArbSetOrGate is
    port (
        clk : in std_logic;
        rst : in std_logic;
        intermediate : in std_logic_vector(1023 downto 0);
        dout : out std_logic
    );
end ArbSetOrGate;


architecture behavioral_ArbSetOrGate of ArbSetOrGate is


signal or_0000_0000 : std_logic := '0';
signal or_0000_0001 : std_logic := '0';
signal or_0000_0002 : std_logic := '0';
signal or_0000_0003 : std_logic := '0';
signal or_0000_0004 : std_logic := '0';
signal or_0000_0005 : std_logic := '0';
signal or_0000_0006 : std_logic := '0';
signal or_0000_0007 : std_logic := '0';
signal or_0000_0008 : std_logic := '0';
signal or_0000_0009 : std_logic := '0';
signal or_0000_0010 : std_logic := '0';
signal or_0000_0011 : std_logic := '0';
signal or_0000_0012 : std_logic := '0';
signal or_0000_0013 : std_logic := '0';
signal or_0000_0014 : std_logic := '0';
signal or_0000_0015 : std_logic := '0';
signal or_0000_0016 : std_logic := '0';
signal or_0000_0017 : std_logic := '0';
signal or_0000_0018 : std_logic := '0';
signal or_0000_0019 : std_logic := '0';
signal or_0000_0020 : std_logic := '0';
signal or_0000_0021 : std_logic := '0';
signal or_0000_0022 : std_logic := '0';
signal or_0000_0023 : std_logic := '0';
signal or_0000_0024 : std_logic := '0';
signal or_0000_0025 : std_logic := '0';
signal or_0000_0026 : std_logic := '0';
signal or_0000_0027 : std_logic := '0';
signal or_0000_0028 : std_logic := '0';
signal or_0000_0029 : std_logic := '0';
signal or_0000_0030 : std_logic := '0';
signal or_0000_0031 : std_logic := '0';
signal or_0000_0032 : std_logic := '0';
signal or_0000_0033 : std_logic := '0';
signal or_0000_0034 : std_logic := '0';
signal or_0000_0035 : std_logic := '0';
signal or_0000_0036 : std_logic := '0';
signal or_0000_0037 : std_logic := '0';
signal or_0000_0038 : std_logic := '0';
signal or_0000_0039 : std_logic := '0';
signal or_0000_0040 : std_logic := '0';
signal or_0000_0041 : std_logic := '0';
signal or_0000_0042 : std_logic := '0';
signal or_0000_0043 : std_logic := '0';
signal or_0000_0044 : std_logic := '0';
signal or_0000_0045 : std_logic := '0';
signal or_0000_0046 : std_logic := '0';
signal or_0000_0047 : std_logic := '0';
signal or_0000_0048 : std_logic := '0';
signal or_0000_0049 : std_logic := '0';
signal or_0000_0050 : std_logic := '0';
signal or_0000_0051 : std_logic := '0';
signal or_0000_0052 : std_logic := '0';
signal or_0000_0053 : std_logic := '0';
signal or_0000_0054 : std_logic := '0';
signal or_0000_0055 : std_logic := '0';
signal or_0000_0056 : std_logic := '0';
signal or_0000_0057 : std_logic := '0';
signal or_0000_0058 : std_logic := '0';
signal or_0000_0059 : std_logic := '0';
signal or_0000_0060 : std_logic := '0';
signal or_0000_0061 : std_logic := '0';
signal or_0000_0062 : std_logic := '0';
signal or_0000_0063 : std_logic := '0';
signal or_0000_0064 : std_logic := '0';
signal or_0000_0065 : std_logic := '0';
signal or_0000_0066 : std_logic := '0';
signal or_0000_0067 : std_logic := '0';
signal or_0000_0068 : std_logic := '0';
signal or_0000_0069 : std_logic := '0';
signal or_0000_0070 : std_logic := '0';
signal or_0000_0071 : std_logic := '0';
signal or_0000_0072 : std_logic := '0';
signal or_0000_0073 : std_logic := '0';
signal or_0000_0074 : std_logic := '0';
signal or_0000_0075 : std_logic := '0';
signal or_0000_0076 : std_logic := '0';
signal or_0000_0077 : std_logic := '0';
signal or_0000_0078 : std_logic := '0';
signal or_0000_0079 : std_logic := '0';
signal or_0000_0080 : std_logic := '0';
signal or_0000_0081 : std_logic := '0';
signal or_0000_0082 : std_logic := '0';
signal or_0000_0083 : std_logic := '0';
signal or_0000_0084 : std_logic := '0';
signal or_0000_0085 : std_logic := '0';
signal or_0000_0086 : std_logic := '0';
signal or_0000_0087 : std_logic := '0';
signal or_0000_0088 : std_logic := '0';
signal or_0000_0089 : std_logic := '0';
signal or_0000_0090 : std_logic := '0';
signal or_0000_0091 : std_logic := '0';
signal or_0000_0092 : std_logic := '0';
signal or_0000_0093 : std_logic := '0';
signal or_0000_0094 : std_logic := '0';
signal or_0000_0095 : std_logic := '0';
signal or_0000_0096 : std_logic := '0';
signal or_0000_0097 : std_logic := '0';
signal or_0000_0098 : std_logic := '0';
signal or_0000_0099 : std_logic := '0';
signal or_0000_0100 : std_logic := '0';
signal or_0000_0101 : std_logic := '0';
signal or_0000_0102 : std_logic := '0';
signal or_0000_0103 : std_logic := '0';
signal or_0000_0104 : std_logic := '0';
signal or_0000_0105 : std_logic := '0';
signal or_0000_0106 : std_logic := '0';
signal or_0000_0107 : std_logic := '0';
signal or_0000_0108 : std_logic := '0';
signal or_0000_0109 : std_logic := '0';
signal or_0000_0110 : std_logic := '0';
signal or_0000_0111 : std_logic := '0';
signal or_0000_0112 : std_logic := '0';
signal or_0000_0113 : std_logic := '0';
signal or_0000_0114 : std_logic := '0';
signal or_0000_0115 : std_logic := '0';
signal or_0000_0116 : std_logic := '0';
signal or_0000_0117 : std_logic := '0';
signal or_0000_0118 : std_logic := '0';
signal or_0000_0119 : std_logic := '0';
signal or_0000_0120 : std_logic := '0';
signal or_0000_0121 : std_logic := '0';
signal or_0000_0122 : std_logic := '0';
signal or_0000_0123 : std_logic := '0';
signal or_0000_0124 : std_logic := '0';
signal or_0000_0125 : std_logic := '0';
signal or_0000_0126 : std_logic := '0';
signal or_0000_0127 : std_logic := '0';
signal or_0000_0128 : std_logic := '0';
signal or_0000_0129 : std_logic := '0';
signal or_0000_0130 : std_logic := '0';
signal or_0000_0131 : std_logic := '0';
signal or_0000_0132 : std_logic := '0';
signal or_0000_0133 : std_logic := '0';
signal or_0000_0134 : std_logic := '0';
signal or_0000_0135 : std_logic := '0';
signal or_0000_0136 : std_logic := '0';
signal or_0000_0137 : std_logic := '0';
signal or_0000_0138 : std_logic := '0';
signal or_0000_0139 : std_logic := '0';
signal or_0000_0140 : std_logic := '0';
signal or_0000_0141 : std_logic := '0';
signal or_0000_0142 : std_logic := '0';
signal or_0000_0143 : std_logic := '0';
signal or_0000_0144 : std_logic := '0';
signal or_0000_0145 : std_logic := '0';
signal or_0000_0146 : std_logic := '0';
signal or_0000_0147 : std_logic := '0';
signal or_0000_0148 : std_logic := '0';
signal or_0000_0149 : std_logic := '0';
signal or_0000_0150 : std_logic := '0';
signal or_0000_0151 : std_logic := '0';
signal or_0000_0152 : std_logic := '0';
signal or_0000_0153 : std_logic := '0';
signal or_0000_0154 : std_logic := '0';
signal or_0000_0155 : std_logic := '0';
signal or_0000_0156 : std_logic := '0';
signal or_0000_0157 : std_logic := '0';
signal or_0000_0158 : std_logic := '0';
signal or_0000_0159 : std_logic := '0';
signal or_0000_0160 : std_logic := '0';
signal or_0000_0161 : std_logic := '0';
signal or_0000_0162 : std_logic := '0';
signal or_0000_0163 : std_logic := '0';
signal or_0000_0164 : std_logic := '0';
signal or_0000_0165 : std_logic := '0';
signal or_0000_0166 : std_logic := '0';
signal or_0000_0167 : std_logic := '0';
signal or_0000_0168 : std_logic := '0';
signal or_0000_0169 : std_logic := '0';
signal or_0000_0170 : std_logic := '0';
signal or_0001_0000 : std_logic := '0';
signal or_0001_0001 : std_logic := '0';
signal or_0001_0002 : std_logic := '0';
signal or_0001_0003 : std_logic := '0';
signal or_0001_0004 : std_logic := '0';
signal or_0001_0005 : std_logic := '0';
signal or_0001_0006 : std_logic := '0';
signal or_0001_0007 : std_logic := '0';
signal or_0001_0008 : std_logic := '0';
signal or_0001_0009 : std_logic := '0';
signal or_0001_0010 : std_logic := '0';
signal or_0001_0011 : std_logic := '0';
signal or_0001_0012 : std_logic := '0';
signal or_0001_0013 : std_logic := '0';
signal or_0001_0014 : std_logic := '0';
signal or_0001_0015 : std_logic := '0';
signal or_0001_0016 : std_logic := '0';
signal or_0001_0017 : std_logic := '0';
signal or_0001_0018 : std_logic := '0';
signal or_0001_0019 : std_logic := '0';
signal or_0001_0020 : std_logic := '0';
signal or_0001_0021 : std_logic := '0';
signal or_0001_0022 : std_logic := '0';
signal or_0001_0023 : std_logic := '0';
signal or_0001_0024 : std_logic := '0';
signal or_0001_0025 : std_logic := '0';
signal or_0001_0026 : std_logic := '0';
signal or_0001_0027 : std_logic := '0';
signal or_0001_0028 : std_logic := '0';
signal or_0002_0000 : std_logic := '0';
signal or_0002_0001 : std_logic := '0';
signal or_0002_0002 : std_logic := '0';
signal or_0002_0003 : std_logic := '0';
signal or_0002_0004 : std_logic := '0';
signal or_0003_0000 : std_logic := '0';


begin


------------------------------------------------------------------------------------------------------------------------
--                                                  RegisteredGates 
------------------------------------------------------------------------------------------------------------------------
INST_or_0000_0000: registeredOR6 port map (clk, rst, intermediate(0), intermediate(1), intermediate(2), intermediate(3), intermediate(4), intermediate(5), or_0000_0000);
INST_or_0000_0001: registeredOR6 port map (clk, rst, intermediate(6), intermediate(7), intermediate(8), intermediate(9), intermediate(10), intermediate(11), or_0000_0001);
INST_or_0000_0002: registeredOR6 port map (clk, rst, intermediate(12), intermediate(13), intermediate(14), intermediate(15), intermediate(16), intermediate(17), or_0000_0002);
INST_or_0000_0003: registeredOR6 port map (clk, rst, intermediate(18), intermediate(19), intermediate(20), intermediate(21), intermediate(22), intermediate(23), or_0000_0003);
INST_or_0000_0004: registeredOR6 port map (clk, rst, intermediate(24), intermediate(25), intermediate(26), intermediate(27), intermediate(28), intermediate(29), or_0000_0004);
INST_or_0000_0005: registeredOR6 port map (clk, rst, intermediate(30), intermediate(31), intermediate(32), intermediate(33), intermediate(34), intermediate(35), or_0000_0005);
INST_or_0000_0006: registeredOR6 port map (clk, rst, intermediate(36), intermediate(37), intermediate(38), intermediate(39), intermediate(40), intermediate(41), or_0000_0006);
INST_or_0000_0007: registeredOR6 port map (clk, rst, intermediate(42), intermediate(43), intermediate(44), intermediate(45), intermediate(46), intermediate(47), or_0000_0007);
INST_or_0000_0008: registeredOR6 port map (clk, rst, intermediate(48), intermediate(49), intermediate(50), intermediate(51), intermediate(52), intermediate(53), or_0000_0008);
INST_or_0000_0009: registeredOR6 port map (clk, rst, intermediate(54), intermediate(55), intermediate(56), intermediate(57), intermediate(58), intermediate(59), or_0000_0009);
INST_or_0000_0010: registeredOR6 port map (clk, rst, intermediate(60), intermediate(61), intermediate(62), intermediate(63), intermediate(64), intermediate(65), or_0000_0010);
INST_or_0000_0011: registeredOR6 port map (clk, rst, intermediate(66), intermediate(67), intermediate(68), intermediate(69), intermediate(70), intermediate(71), or_0000_0011);
INST_or_0000_0012: registeredOR6 port map (clk, rst, intermediate(72), intermediate(73), intermediate(74), intermediate(75), intermediate(76), intermediate(77), or_0000_0012);
INST_or_0000_0013: registeredOR6 port map (clk, rst, intermediate(78), intermediate(79), intermediate(80), intermediate(81), intermediate(82), intermediate(83), or_0000_0013);
INST_or_0000_0014: registeredOR6 port map (clk, rst, intermediate(84), intermediate(85), intermediate(86), intermediate(87), intermediate(88), intermediate(89), or_0000_0014);
INST_or_0000_0015: registeredOR6 port map (clk, rst, intermediate(90), intermediate(91), intermediate(92), intermediate(93), intermediate(94), intermediate(95), or_0000_0015);
INST_or_0000_0016: registeredOR6 port map (clk, rst, intermediate(96), intermediate(97), intermediate(98), intermediate(99), intermediate(100), intermediate(101), or_0000_0016);
INST_or_0000_0017: registeredOR6 port map (clk, rst, intermediate(102), intermediate(103), intermediate(104), intermediate(105), intermediate(106), intermediate(107), or_0000_0017);
INST_or_0000_0018: registeredOR6 port map (clk, rst, intermediate(108), intermediate(109), intermediate(110), intermediate(111), intermediate(112), intermediate(113), or_0000_0018);
INST_or_0000_0019: registeredOR6 port map (clk, rst, intermediate(114), intermediate(115), intermediate(116), intermediate(117), intermediate(118), intermediate(119), or_0000_0019);
INST_or_0000_0020: registeredOR6 port map (clk, rst, intermediate(120), intermediate(121), intermediate(122), intermediate(123), intermediate(124), intermediate(125), or_0000_0020);
INST_or_0000_0021: registeredOR6 port map (clk, rst, intermediate(126), intermediate(127), intermediate(128), intermediate(129), intermediate(130), intermediate(131), or_0000_0021);
INST_or_0000_0022: registeredOR6 port map (clk, rst, intermediate(132), intermediate(133), intermediate(134), intermediate(135), intermediate(136), intermediate(137), or_0000_0022);
INST_or_0000_0023: registeredOR6 port map (clk, rst, intermediate(138), intermediate(139), intermediate(140), intermediate(141), intermediate(142), intermediate(143), or_0000_0023);
INST_or_0000_0024: registeredOR6 port map (clk, rst, intermediate(144), intermediate(145), intermediate(146), intermediate(147), intermediate(148), intermediate(149), or_0000_0024);
INST_or_0000_0025: registeredOR6 port map (clk, rst, intermediate(150), intermediate(151), intermediate(152), intermediate(153), intermediate(154), intermediate(155), or_0000_0025);
INST_or_0000_0026: registeredOR6 port map (clk, rst, intermediate(156), intermediate(157), intermediate(158), intermediate(159), intermediate(160), intermediate(161), or_0000_0026);
INST_or_0000_0027: registeredOR6 port map (clk, rst, intermediate(162), intermediate(163), intermediate(164), intermediate(165), intermediate(166), intermediate(167), or_0000_0027);
INST_or_0000_0028: registeredOR6 port map (clk, rst, intermediate(168), intermediate(169), intermediate(170), intermediate(171), intermediate(172), intermediate(173), or_0000_0028);
INST_or_0000_0029: registeredOR6 port map (clk, rst, intermediate(174), intermediate(175), intermediate(176), intermediate(177), intermediate(178), intermediate(179), or_0000_0029);
INST_or_0000_0030: registeredOR6 port map (clk, rst, intermediate(180), intermediate(181), intermediate(182), intermediate(183), intermediate(184), intermediate(185), or_0000_0030);
INST_or_0000_0031: registeredOR6 port map (clk, rst, intermediate(186), intermediate(187), intermediate(188), intermediate(189), intermediate(190), intermediate(191), or_0000_0031);
INST_or_0000_0032: registeredOR6 port map (clk, rst, intermediate(192), intermediate(193), intermediate(194), intermediate(195), intermediate(196), intermediate(197), or_0000_0032);
INST_or_0000_0033: registeredOR6 port map (clk, rst, intermediate(198), intermediate(199), intermediate(200), intermediate(201), intermediate(202), intermediate(203), or_0000_0033);
INST_or_0000_0034: registeredOR6 port map (clk, rst, intermediate(204), intermediate(205), intermediate(206), intermediate(207), intermediate(208), intermediate(209), or_0000_0034);
INST_or_0000_0035: registeredOR6 port map (clk, rst, intermediate(210), intermediate(211), intermediate(212), intermediate(213), intermediate(214), intermediate(215), or_0000_0035);
INST_or_0000_0036: registeredOR6 port map (clk, rst, intermediate(216), intermediate(217), intermediate(218), intermediate(219), intermediate(220), intermediate(221), or_0000_0036);
INST_or_0000_0037: registeredOR6 port map (clk, rst, intermediate(222), intermediate(223), intermediate(224), intermediate(225), intermediate(226), intermediate(227), or_0000_0037);
INST_or_0000_0038: registeredOR6 port map (clk, rst, intermediate(228), intermediate(229), intermediate(230), intermediate(231), intermediate(232), intermediate(233), or_0000_0038);
INST_or_0000_0039: registeredOR6 port map (clk, rst, intermediate(234), intermediate(235), intermediate(236), intermediate(237), intermediate(238), intermediate(239), or_0000_0039);
INST_or_0000_0040: registeredOR6 port map (clk, rst, intermediate(240), intermediate(241), intermediate(242), intermediate(243), intermediate(244), intermediate(245), or_0000_0040);
INST_or_0000_0041: registeredOR6 port map (clk, rst, intermediate(246), intermediate(247), intermediate(248), intermediate(249), intermediate(250), intermediate(251), or_0000_0041);
INST_or_0000_0042: registeredOR6 port map (clk, rst, intermediate(252), intermediate(253), intermediate(254), intermediate(255), intermediate(256), intermediate(257), or_0000_0042);
INST_or_0000_0043: registeredOR6 port map (clk, rst, intermediate(258), intermediate(259), intermediate(260), intermediate(261), intermediate(262), intermediate(263), or_0000_0043);
INST_or_0000_0044: registeredOR6 port map (clk, rst, intermediate(264), intermediate(265), intermediate(266), intermediate(267), intermediate(268), intermediate(269), or_0000_0044);
INST_or_0000_0045: registeredOR6 port map (clk, rst, intermediate(270), intermediate(271), intermediate(272), intermediate(273), intermediate(274), intermediate(275), or_0000_0045);
INST_or_0000_0046: registeredOR6 port map (clk, rst, intermediate(276), intermediate(277), intermediate(278), intermediate(279), intermediate(280), intermediate(281), or_0000_0046);
INST_or_0000_0047: registeredOR6 port map (clk, rst, intermediate(282), intermediate(283), intermediate(284), intermediate(285), intermediate(286), intermediate(287), or_0000_0047);
INST_or_0000_0048: registeredOR6 port map (clk, rst, intermediate(288), intermediate(289), intermediate(290), intermediate(291), intermediate(292), intermediate(293), or_0000_0048);
INST_or_0000_0049: registeredOR6 port map (clk, rst, intermediate(294), intermediate(295), intermediate(296), intermediate(297), intermediate(298), intermediate(299), or_0000_0049);
INST_or_0000_0050: registeredOR6 port map (clk, rst, intermediate(300), intermediate(301), intermediate(302), intermediate(303), intermediate(304), intermediate(305), or_0000_0050);
INST_or_0000_0051: registeredOR6 port map (clk, rst, intermediate(306), intermediate(307), intermediate(308), intermediate(309), intermediate(310), intermediate(311), or_0000_0051);
INST_or_0000_0052: registeredOR6 port map (clk, rst, intermediate(312), intermediate(313), intermediate(314), intermediate(315), intermediate(316), intermediate(317), or_0000_0052);
INST_or_0000_0053: registeredOR6 port map (clk, rst, intermediate(318), intermediate(319), intermediate(320), intermediate(321), intermediate(322), intermediate(323), or_0000_0053);
INST_or_0000_0054: registeredOR6 port map (clk, rst, intermediate(324), intermediate(325), intermediate(326), intermediate(327), intermediate(328), intermediate(329), or_0000_0054);
INST_or_0000_0055: registeredOR6 port map (clk, rst, intermediate(330), intermediate(331), intermediate(332), intermediate(333), intermediate(334), intermediate(335), or_0000_0055);
INST_or_0000_0056: registeredOR6 port map (clk, rst, intermediate(336), intermediate(337), intermediate(338), intermediate(339), intermediate(340), intermediate(341), or_0000_0056);
INST_or_0000_0057: registeredOR6 port map (clk, rst, intermediate(342), intermediate(343), intermediate(344), intermediate(345), intermediate(346), intermediate(347), or_0000_0057);
INST_or_0000_0058: registeredOR6 port map (clk, rst, intermediate(348), intermediate(349), intermediate(350), intermediate(351), intermediate(352), intermediate(353), or_0000_0058);
INST_or_0000_0059: registeredOR6 port map (clk, rst, intermediate(354), intermediate(355), intermediate(356), intermediate(357), intermediate(358), intermediate(359), or_0000_0059);
INST_or_0000_0060: registeredOR6 port map (clk, rst, intermediate(360), intermediate(361), intermediate(362), intermediate(363), intermediate(364), intermediate(365), or_0000_0060);
INST_or_0000_0061: registeredOR6 port map (clk, rst, intermediate(366), intermediate(367), intermediate(368), intermediate(369), intermediate(370), intermediate(371), or_0000_0061);
INST_or_0000_0062: registeredOR6 port map (clk, rst, intermediate(372), intermediate(373), intermediate(374), intermediate(375), intermediate(376), intermediate(377), or_0000_0062);
INST_or_0000_0063: registeredOR6 port map (clk, rst, intermediate(378), intermediate(379), intermediate(380), intermediate(381), intermediate(382), intermediate(383), or_0000_0063);
INST_or_0000_0064: registeredOR6 port map (clk, rst, intermediate(384), intermediate(385), intermediate(386), intermediate(387), intermediate(388), intermediate(389), or_0000_0064);
INST_or_0000_0065: registeredOR6 port map (clk, rst, intermediate(390), intermediate(391), intermediate(392), intermediate(393), intermediate(394), intermediate(395), or_0000_0065);
INST_or_0000_0066: registeredOR6 port map (clk, rst, intermediate(396), intermediate(397), intermediate(398), intermediate(399), intermediate(400), intermediate(401), or_0000_0066);
INST_or_0000_0067: registeredOR6 port map (clk, rst, intermediate(402), intermediate(403), intermediate(404), intermediate(405), intermediate(406), intermediate(407), or_0000_0067);
INST_or_0000_0068: registeredOR6 port map (clk, rst, intermediate(408), intermediate(409), intermediate(410), intermediate(411), intermediate(412), intermediate(413), or_0000_0068);
INST_or_0000_0069: registeredOR6 port map (clk, rst, intermediate(414), intermediate(415), intermediate(416), intermediate(417), intermediate(418), intermediate(419), or_0000_0069);
INST_or_0000_0070: registeredOR6 port map (clk, rst, intermediate(420), intermediate(421), intermediate(422), intermediate(423), intermediate(424), intermediate(425), or_0000_0070);
INST_or_0000_0071: registeredOR6 port map (clk, rst, intermediate(426), intermediate(427), intermediate(428), intermediate(429), intermediate(430), intermediate(431), or_0000_0071);
INST_or_0000_0072: registeredOR6 port map (clk, rst, intermediate(432), intermediate(433), intermediate(434), intermediate(435), intermediate(436), intermediate(437), or_0000_0072);
INST_or_0000_0073: registeredOR6 port map (clk, rst, intermediate(438), intermediate(439), intermediate(440), intermediate(441), intermediate(442), intermediate(443), or_0000_0073);
INST_or_0000_0074: registeredOR6 port map (clk, rst, intermediate(444), intermediate(445), intermediate(446), intermediate(447), intermediate(448), intermediate(449), or_0000_0074);
INST_or_0000_0075: registeredOR6 port map (clk, rst, intermediate(450), intermediate(451), intermediate(452), intermediate(453), intermediate(454), intermediate(455), or_0000_0075);
INST_or_0000_0076: registeredOR6 port map (clk, rst, intermediate(456), intermediate(457), intermediate(458), intermediate(459), intermediate(460), intermediate(461), or_0000_0076);
INST_or_0000_0077: registeredOR6 port map (clk, rst, intermediate(462), intermediate(463), intermediate(464), intermediate(465), intermediate(466), intermediate(467), or_0000_0077);
INST_or_0000_0078: registeredOR6 port map (clk, rst, intermediate(468), intermediate(469), intermediate(470), intermediate(471), intermediate(472), intermediate(473), or_0000_0078);
INST_or_0000_0079: registeredOR6 port map (clk, rst, intermediate(474), intermediate(475), intermediate(476), intermediate(477), intermediate(478), intermediate(479), or_0000_0079);
INST_or_0000_0080: registeredOR6 port map (clk, rst, intermediate(480), intermediate(481), intermediate(482), intermediate(483), intermediate(484), intermediate(485), or_0000_0080);
INST_or_0000_0081: registeredOR6 port map (clk, rst, intermediate(486), intermediate(487), intermediate(488), intermediate(489), intermediate(490), intermediate(491), or_0000_0081);
INST_or_0000_0082: registeredOR6 port map (clk, rst, intermediate(492), intermediate(493), intermediate(494), intermediate(495), intermediate(496), intermediate(497), or_0000_0082);
INST_or_0000_0083: registeredOR6 port map (clk, rst, intermediate(498), intermediate(499), intermediate(500), intermediate(501), intermediate(502), intermediate(503), or_0000_0083);
INST_or_0000_0084: registeredOR6 port map (clk, rst, intermediate(504), intermediate(505), intermediate(506), intermediate(507), intermediate(508), intermediate(509), or_0000_0084);
INST_or_0000_0085: registeredOR6 port map (clk, rst, intermediate(510), intermediate(511), intermediate(512), intermediate(513), intermediate(514), intermediate(515), or_0000_0085);
INST_or_0000_0086: registeredOR6 port map (clk, rst, intermediate(516), intermediate(517), intermediate(518), intermediate(519), intermediate(520), intermediate(521), or_0000_0086);
INST_or_0000_0087: registeredOR6 port map (clk, rst, intermediate(522), intermediate(523), intermediate(524), intermediate(525), intermediate(526), intermediate(527), or_0000_0087);
INST_or_0000_0088: registeredOR6 port map (clk, rst, intermediate(528), intermediate(529), intermediate(530), intermediate(531), intermediate(532), intermediate(533), or_0000_0088);
INST_or_0000_0089: registeredOR6 port map (clk, rst, intermediate(534), intermediate(535), intermediate(536), intermediate(537), intermediate(538), intermediate(539), or_0000_0089);
INST_or_0000_0090: registeredOR6 port map (clk, rst, intermediate(540), intermediate(541), intermediate(542), intermediate(543), intermediate(544), intermediate(545), or_0000_0090);
INST_or_0000_0091: registeredOR6 port map (clk, rst, intermediate(546), intermediate(547), intermediate(548), intermediate(549), intermediate(550), intermediate(551), or_0000_0091);
INST_or_0000_0092: registeredOR6 port map (clk, rst, intermediate(552), intermediate(553), intermediate(554), intermediate(555), intermediate(556), intermediate(557), or_0000_0092);
INST_or_0000_0093: registeredOR6 port map (clk, rst, intermediate(558), intermediate(559), intermediate(560), intermediate(561), intermediate(562), intermediate(563), or_0000_0093);
INST_or_0000_0094: registeredOR6 port map (clk, rst, intermediate(564), intermediate(565), intermediate(566), intermediate(567), intermediate(568), intermediate(569), or_0000_0094);
INST_or_0000_0095: registeredOR6 port map (clk, rst, intermediate(570), intermediate(571), intermediate(572), intermediate(573), intermediate(574), intermediate(575), or_0000_0095);
INST_or_0000_0096: registeredOR6 port map (clk, rst, intermediate(576), intermediate(577), intermediate(578), intermediate(579), intermediate(580), intermediate(581), or_0000_0096);
INST_or_0000_0097: registeredOR6 port map (clk, rst, intermediate(582), intermediate(583), intermediate(584), intermediate(585), intermediate(586), intermediate(587), or_0000_0097);
INST_or_0000_0098: registeredOR6 port map (clk, rst, intermediate(588), intermediate(589), intermediate(590), intermediate(591), intermediate(592), intermediate(593), or_0000_0098);
INST_or_0000_0099: registeredOR6 port map (clk, rst, intermediate(594), intermediate(595), intermediate(596), intermediate(597), intermediate(598), intermediate(599), or_0000_0099);
INST_or_0000_0100: registeredOR6 port map (clk, rst, intermediate(600), intermediate(601), intermediate(602), intermediate(603), intermediate(604), intermediate(605), or_0000_0100);
INST_or_0000_0101: registeredOR6 port map (clk, rst, intermediate(606), intermediate(607), intermediate(608), intermediate(609), intermediate(610), intermediate(611), or_0000_0101);
INST_or_0000_0102: registeredOR6 port map (clk, rst, intermediate(612), intermediate(613), intermediate(614), intermediate(615), intermediate(616), intermediate(617), or_0000_0102);
INST_or_0000_0103: registeredOR6 port map (clk, rst, intermediate(618), intermediate(619), intermediate(620), intermediate(621), intermediate(622), intermediate(623), or_0000_0103);
INST_or_0000_0104: registeredOR6 port map (clk, rst, intermediate(624), intermediate(625), intermediate(626), intermediate(627), intermediate(628), intermediate(629), or_0000_0104);
INST_or_0000_0105: registeredOR6 port map (clk, rst, intermediate(630), intermediate(631), intermediate(632), intermediate(633), intermediate(634), intermediate(635), or_0000_0105);
INST_or_0000_0106: registeredOR6 port map (clk, rst, intermediate(636), intermediate(637), intermediate(638), intermediate(639), intermediate(640), intermediate(641), or_0000_0106);
INST_or_0000_0107: registeredOR6 port map (clk, rst, intermediate(642), intermediate(643), intermediate(644), intermediate(645), intermediate(646), intermediate(647), or_0000_0107);
INST_or_0000_0108: registeredOR6 port map (clk, rst, intermediate(648), intermediate(649), intermediate(650), intermediate(651), intermediate(652), intermediate(653), or_0000_0108);
INST_or_0000_0109: registeredOR6 port map (clk, rst, intermediate(654), intermediate(655), intermediate(656), intermediate(657), intermediate(658), intermediate(659), or_0000_0109);
INST_or_0000_0110: registeredOR6 port map (clk, rst, intermediate(660), intermediate(661), intermediate(662), intermediate(663), intermediate(664), intermediate(665), or_0000_0110);
INST_or_0000_0111: registeredOR6 port map (clk, rst, intermediate(666), intermediate(667), intermediate(668), intermediate(669), intermediate(670), intermediate(671), or_0000_0111);
INST_or_0000_0112: registeredOR6 port map (clk, rst, intermediate(672), intermediate(673), intermediate(674), intermediate(675), intermediate(676), intermediate(677), or_0000_0112);
INST_or_0000_0113: registeredOR6 port map (clk, rst, intermediate(678), intermediate(679), intermediate(680), intermediate(681), intermediate(682), intermediate(683), or_0000_0113);
INST_or_0000_0114: registeredOR6 port map (clk, rst, intermediate(684), intermediate(685), intermediate(686), intermediate(687), intermediate(688), intermediate(689), or_0000_0114);
INST_or_0000_0115: registeredOR6 port map (clk, rst, intermediate(690), intermediate(691), intermediate(692), intermediate(693), intermediate(694), intermediate(695), or_0000_0115);
INST_or_0000_0116: registeredOR6 port map (clk, rst, intermediate(696), intermediate(697), intermediate(698), intermediate(699), intermediate(700), intermediate(701), or_0000_0116);
INST_or_0000_0117: registeredOR6 port map (clk, rst, intermediate(702), intermediate(703), intermediate(704), intermediate(705), intermediate(706), intermediate(707), or_0000_0117);
INST_or_0000_0118: registeredOR6 port map (clk, rst, intermediate(708), intermediate(709), intermediate(710), intermediate(711), intermediate(712), intermediate(713), or_0000_0118);
INST_or_0000_0119: registeredOR6 port map (clk, rst, intermediate(714), intermediate(715), intermediate(716), intermediate(717), intermediate(718), intermediate(719), or_0000_0119);
INST_or_0000_0120: registeredOR6 port map (clk, rst, intermediate(720), intermediate(721), intermediate(722), intermediate(723), intermediate(724), intermediate(725), or_0000_0120);
INST_or_0000_0121: registeredOR6 port map (clk, rst, intermediate(726), intermediate(727), intermediate(728), intermediate(729), intermediate(730), intermediate(731), or_0000_0121);
INST_or_0000_0122: registeredOR6 port map (clk, rst, intermediate(732), intermediate(733), intermediate(734), intermediate(735), intermediate(736), intermediate(737), or_0000_0122);
INST_or_0000_0123: registeredOR6 port map (clk, rst, intermediate(738), intermediate(739), intermediate(740), intermediate(741), intermediate(742), intermediate(743), or_0000_0123);
INST_or_0000_0124: registeredOR6 port map (clk, rst, intermediate(744), intermediate(745), intermediate(746), intermediate(747), intermediate(748), intermediate(749), or_0000_0124);
INST_or_0000_0125: registeredOR6 port map (clk, rst, intermediate(750), intermediate(751), intermediate(752), intermediate(753), intermediate(754), intermediate(755), or_0000_0125);
INST_or_0000_0126: registeredOR6 port map (clk, rst, intermediate(756), intermediate(757), intermediate(758), intermediate(759), intermediate(760), intermediate(761), or_0000_0126);
INST_or_0000_0127: registeredOR6 port map (clk, rst, intermediate(762), intermediate(763), intermediate(764), intermediate(765), intermediate(766), intermediate(767), or_0000_0127);
INST_or_0000_0128: registeredOR6 port map (clk, rst, intermediate(768), intermediate(769), intermediate(770), intermediate(771), intermediate(772), intermediate(773), or_0000_0128);
INST_or_0000_0129: registeredOR6 port map (clk, rst, intermediate(774), intermediate(775), intermediate(776), intermediate(777), intermediate(778), intermediate(779), or_0000_0129);
INST_or_0000_0130: registeredOR6 port map (clk, rst, intermediate(780), intermediate(781), intermediate(782), intermediate(783), intermediate(784), intermediate(785), or_0000_0130);
INST_or_0000_0131: registeredOR6 port map (clk, rst, intermediate(786), intermediate(787), intermediate(788), intermediate(789), intermediate(790), intermediate(791), or_0000_0131);
INST_or_0000_0132: registeredOR6 port map (clk, rst, intermediate(792), intermediate(793), intermediate(794), intermediate(795), intermediate(796), intermediate(797), or_0000_0132);
INST_or_0000_0133: registeredOR6 port map (clk, rst, intermediate(798), intermediate(799), intermediate(800), intermediate(801), intermediate(802), intermediate(803), or_0000_0133);
INST_or_0000_0134: registeredOR6 port map (clk, rst, intermediate(804), intermediate(805), intermediate(806), intermediate(807), intermediate(808), intermediate(809), or_0000_0134);
INST_or_0000_0135: registeredOR6 port map (clk, rst, intermediate(810), intermediate(811), intermediate(812), intermediate(813), intermediate(814), intermediate(815), or_0000_0135);
INST_or_0000_0136: registeredOR6 port map (clk, rst, intermediate(816), intermediate(817), intermediate(818), intermediate(819), intermediate(820), intermediate(821), or_0000_0136);
INST_or_0000_0137: registeredOR6 port map (clk, rst, intermediate(822), intermediate(823), intermediate(824), intermediate(825), intermediate(826), intermediate(827), or_0000_0137);
INST_or_0000_0138: registeredOR6 port map (clk, rst, intermediate(828), intermediate(829), intermediate(830), intermediate(831), intermediate(832), intermediate(833), or_0000_0138);
INST_or_0000_0139: registeredOR6 port map (clk, rst, intermediate(834), intermediate(835), intermediate(836), intermediate(837), intermediate(838), intermediate(839), or_0000_0139);
INST_or_0000_0140: registeredOR6 port map (clk, rst, intermediate(840), intermediate(841), intermediate(842), intermediate(843), intermediate(844), intermediate(845), or_0000_0140);
INST_or_0000_0141: registeredOR6 port map (clk, rst, intermediate(846), intermediate(847), intermediate(848), intermediate(849), intermediate(850), intermediate(851), or_0000_0141);
INST_or_0000_0142: registeredOR6 port map (clk, rst, intermediate(852), intermediate(853), intermediate(854), intermediate(855), intermediate(856), intermediate(857), or_0000_0142);
INST_or_0000_0143: registeredOR6 port map (clk, rst, intermediate(858), intermediate(859), intermediate(860), intermediate(861), intermediate(862), intermediate(863), or_0000_0143);
INST_or_0000_0144: registeredOR6 port map (clk, rst, intermediate(864), intermediate(865), intermediate(866), intermediate(867), intermediate(868), intermediate(869), or_0000_0144);
INST_or_0000_0145: registeredOR6 port map (clk, rst, intermediate(870), intermediate(871), intermediate(872), intermediate(873), intermediate(874), intermediate(875), or_0000_0145);
INST_or_0000_0146: registeredOR6 port map (clk, rst, intermediate(876), intermediate(877), intermediate(878), intermediate(879), intermediate(880), intermediate(881), or_0000_0146);
INST_or_0000_0147: registeredOR6 port map (clk, rst, intermediate(882), intermediate(883), intermediate(884), intermediate(885), intermediate(886), intermediate(887), or_0000_0147);
INST_or_0000_0148: registeredOR6 port map (clk, rst, intermediate(888), intermediate(889), intermediate(890), intermediate(891), intermediate(892), intermediate(893), or_0000_0148);
INST_or_0000_0149: registeredOR6 port map (clk, rst, intermediate(894), intermediate(895), intermediate(896), intermediate(897), intermediate(898), intermediate(899), or_0000_0149);
INST_or_0000_0150: registeredOR6 port map (clk, rst, intermediate(900), intermediate(901), intermediate(902), intermediate(903), intermediate(904), intermediate(905), or_0000_0150);
INST_or_0000_0151: registeredOR6 port map (clk, rst, intermediate(906), intermediate(907), intermediate(908), intermediate(909), intermediate(910), intermediate(911), or_0000_0151);
INST_or_0000_0152: registeredOR6 port map (clk, rst, intermediate(912), intermediate(913), intermediate(914), intermediate(915), intermediate(916), intermediate(917), or_0000_0152);
INST_or_0000_0153: registeredOR6 port map (clk, rst, intermediate(918), intermediate(919), intermediate(920), intermediate(921), intermediate(922), intermediate(923), or_0000_0153);
INST_or_0000_0154: registeredOR6 port map (clk, rst, intermediate(924), intermediate(925), intermediate(926), intermediate(927), intermediate(928), intermediate(929), or_0000_0154);
INST_or_0000_0155: registeredOR6 port map (clk, rst, intermediate(930), intermediate(931), intermediate(932), intermediate(933), intermediate(934), intermediate(935), or_0000_0155);
INST_or_0000_0156: registeredOR6 port map (clk, rst, intermediate(936), intermediate(937), intermediate(938), intermediate(939), intermediate(940), intermediate(941), or_0000_0156);
INST_or_0000_0157: registeredOR6 port map (clk, rst, intermediate(942), intermediate(943), intermediate(944), intermediate(945), intermediate(946), intermediate(947), or_0000_0157);
INST_or_0000_0158: registeredOR6 port map (clk, rst, intermediate(948), intermediate(949), intermediate(950), intermediate(951), intermediate(952), intermediate(953), or_0000_0158);
INST_or_0000_0159: registeredOR6 port map (clk, rst, intermediate(954), intermediate(955), intermediate(956), intermediate(957), intermediate(958), intermediate(959), or_0000_0159);
INST_or_0000_0160: registeredOR6 port map (clk, rst, intermediate(960), intermediate(961), intermediate(962), intermediate(963), intermediate(964), intermediate(965), or_0000_0160);
INST_or_0000_0161: registeredOR6 port map (clk, rst, intermediate(966), intermediate(967), intermediate(968), intermediate(969), intermediate(970), intermediate(971), or_0000_0161);
INST_or_0000_0162: registeredOR6 port map (clk, rst, intermediate(972), intermediate(973), intermediate(974), intermediate(975), intermediate(976), intermediate(977), or_0000_0162);
INST_or_0000_0163: registeredOR6 port map (clk, rst, intermediate(978), intermediate(979), intermediate(980), intermediate(981), intermediate(982), intermediate(983), or_0000_0163);
INST_or_0000_0164: registeredOR6 port map (clk, rst, intermediate(984), intermediate(985), intermediate(986), intermediate(987), intermediate(988), intermediate(989), or_0000_0164);
INST_or_0000_0165: registeredOR6 port map (clk, rst, intermediate(990), intermediate(991), intermediate(992), intermediate(993), intermediate(994), intermediate(995), or_0000_0165);
INST_or_0000_0166: registeredOR6 port map (clk, rst, intermediate(996), intermediate(997), intermediate(998), intermediate(999), intermediate(1000), intermediate(1001), or_0000_0166);
INST_or_0000_0167: registeredOR6 port map (clk, rst, intermediate(1002), intermediate(1003), intermediate(1004), intermediate(1005), intermediate(1006), intermediate(1007), or_0000_0167);
INST_or_0000_0168: registeredOR6 port map (clk, rst, intermediate(1008), intermediate(1009), intermediate(1010), intermediate(1011), intermediate(1012), intermediate(1013), or_0000_0168);
INST_or_0000_0169: registeredOR6 port map (clk, rst, intermediate(1014), intermediate(1015), intermediate(1016), intermediate(1017), intermediate(1018), intermediate(1019), or_0000_0169);
INST_or_0000_0170: registeredOR4 port map (clk, rst, intermediate(1020), intermediate(1021), intermediate(1022), intermediate(1023), or_0000_0170);
INST_or_0001_0000: registeredOR6 port map (clk, rst, or_0000_0000, or_0000_0001, or_0000_0002, or_0000_0003, or_0000_0004, or_0000_0005, or_0001_0000);
INST_or_0001_0001: registeredOR6 port map (clk, rst, or_0000_0006, or_0000_0007, or_0000_0008, or_0000_0009, or_0000_0010, or_0000_0011, or_0001_0001);
INST_or_0001_0002: registeredOR6 port map (clk, rst, or_0000_0012, or_0000_0013, or_0000_0014, or_0000_0015, or_0000_0016, or_0000_0017, or_0001_0002);
INST_or_0001_0003: registeredOR6 port map (clk, rst, or_0000_0018, or_0000_0019, or_0000_0020, or_0000_0021, or_0000_0022, or_0000_0023, or_0001_0003);
INST_or_0001_0004: registeredOR6 port map (clk, rst, or_0000_0024, or_0000_0025, or_0000_0026, or_0000_0027, or_0000_0028, or_0000_0029, or_0001_0004);
INST_or_0001_0005: registeredOR6 port map (clk, rst, or_0000_0030, or_0000_0031, or_0000_0032, or_0000_0033, or_0000_0034, or_0000_0035, or_0001_0005);
INST_or_0001_0006: registeredOR6 port map (clk, rst, or_0000_0036, or_0000_0037, or_0000_0038, or_0000_0039, or_0000_0040, or_0000_0041, or_0001_0006);
INST_or_0001_0007: registeredOR6 port map (clk, rst, or_0000_0042, or_0000_0043, or_0000_0044, or_0000_0045, or_0000_0046, or_0000_0047, or_0001_0007);
INST_or_0001_0008: registeredOR6 port map (clk, rst, or_0000_0048, or_0000_0049, or_0000_0050, or_0000_0051, or_0000_0052, or_0000_0053, or_0001_0008);
INST_or_0001_0009: registeredOR6 port map (clk, rst, or_0000_0054, or_0000_0055, or_0000_0056, or_0000_0057, or_0000_0058, or_0000_0059, or_0001_0009);
INST_or_0001_0010: registeredOR6 port map (clk, rst, or_0000_0060, or_0000_0061, or_0000_0062, or_0000_0063, or_0000_0064, or_0000_0065, or_0001_0010);
INST_or_0001_0011: registeredOR6 port map (clk, rst, or_0000_0066, or_0000_0067, or_0000_0068, or_0000_0069, or_0000_0070, or_0000_0071, or_0001_0011);
INST_or_0001_0012: registeredOR6 port map (clk, rst, or_0000_0072, or_0000_0073, or_0000_0074, or_0000_0075, or_0000_0076, or_0000_0077, or_0001_0012);
INST_or_0001_0013: registeredOR6 port map (clk, rst, or_0000_0078, or_0000_0079, or_0000_0080, or_0000_0081, or_0000_0082, or_0000_0083, or_0001_0013);
INST_or_0001_0014: registeredOR6 port map (clk, rst, or_0000_0084, or_0000_0085, or_0000_0086, or_0000_0087, or_0000_0088, or_0000_0089, or_0001_0014);
INST_or_0001_0015: registeredOR6 port map (clk, rst, or_0000_0090, or_0000_0091, or_0000_0092, or_0000_0093, or_0000_0094, or_0000_0095, or_0001_0015);
INST_or_0001_0016: registeredOR6 port map (clk, rst, or_0000_0096, or_0000_0097, or_0000_0098, or_0000_0099, or_0000_0100, or_0000_0101, or_0001_0016);
INST_or_0001_0017: registeredOR6 port map (clk, rst, or_0000_0102, or_0000_0103, or_0000_0104, or_0000_0105, or_0000_0106, or_0000_0107, or_0001_0017);
INST_or_0001_0018: registeredOR6 port map (clk, rst, or_0000_0108, or_0000_0109, or_0000_0110, or_0000_0111, or_0000_0112, or_0000_0113, or_0001_0018);
INST_or_0001_0019: registeredOR6 port map (clk, rst, or_0000_0114, or_0000_0115, or_0000_0116, or_0000_0117, or_0000_0118, or_0000_0119, or_0001_0019);
INST_or_0001_0020: registeredOR6 port map (clk, rst, or_0000_0120, or_0000_0121, or_0000_0122, or_0000_0123, or_0000_0124, or_0000_0125, or_0001_0020);
INST_or_0001_0021: registeredOR6 port map (clk, rst, or_0000_0126, or_0000_0127, or_0000_0128, or_0000_0129, or_0000_0130, or_0000_0131, or_0001_0021);
INST_or_0001_0022: registeredOR6 port map (clk, rst, or_0000_0132, or_0000_0133, or_0000_0134, or_0000_0135, or_0000_0136, or_0000_0137, or_0001_0022);
INST_or_0001_0023: registeredOR6 port map (clk, rst, or_0000_0138, or_0000_0139, or_0000_0140, or_0000_0141, or_0000_0142, or_0000_0143, or_0001_0023);
INST_or_0001_0024: registeredOR6 port map (clk, rst, or_0000_0144, or_0000_0145, or_0000_0146, or_0000_0147, or_0000_0148, or_0000_0149, or_0001_0024);
INST_or_0001_0025: registeredOR6 port map (clk, rst, or_0000_0150, or_0000_0151, or_0000_0152, or_0000_0153, or_0000_0154, or_0000_0155, or_0001_0025);
INST_or_0001_0026: registeredOR6 port map (clk, rst, or_0000_0156, or_0000_0157, or_0000_0158, or_0000_0159, or_0000_0160, or_0000_0161, or_0001_0026);
INST_or_0001_0027: registeredOR6 port map (clk, rst, or_0000_0162, or_0000_0163, or_0000_0164, or_0000_0165, or_0000_0166, or_0000_0167, or_0001_0027);
INST_or_0001_0028: registeredOR3 port map (clk, rst, or_0000_0168, or_0000_0169, or_0000_0170, or_0001_0028);
INST_or_0002_0000: registeredOR6 port map (clk, rst, or_0001_0000, or_0001_0001, or_0001_0002, or_0001_0003, or_0001_0004, or_0001_0005, or_0002_0000);
INST_or_0002_0001: registeredOR6 port map (clk, rst, or_0001_0006, or_0001_0007, or_0001_0008, or_0001_0009, or_0001_0010, or_0001_0011, or_0002_0001);
INST_or_0002_0002: registeredOR6 port map (clk, rst, or_0001_0012, or_0001_0013, or_0001_0014, or_0001_0015, or_0001_0016, or_0001_0017, or_0002_0002);
INST_or_0002_0003: registeredOR6 port map (clk, rst, or_0001_0018, or_0001_0019, or_0001_0020, or_0001_0021, or_0001_0022, or_0001_0023, or_0002_0003);
INST_or_0002_0004: registeredOR5 port map (clk, rst, or_0001_0024, or_0001_0025, or_0001_0026, or_0001_0027, or_0001_0028, or_0002_0004);
INST_or_0003_0000: registeredOR5 port map (clk, rst, or_0002_0000, or_0002_0001, or_0002_0002, or_0002_0003, or_0002_0004, or_0003_0000);

------------------------------------------------------------------------------------------------------------------------
--                                                   Drive Outputs 
------------------------------------------------------------------------------------------------------------------------
dout <= or_0003_0000;

end behavioral_ArbSetOrGate;

