library IEEE;
use IEEE.std_logic_1164.ALL;
use IEEE.numeric_std.ALL;


entity CrossClockStdLogic is
    port (
        clk : in std_logic;
        rst : in std_logic
    );
end CrossClockStdLogic;


architecture behavioral_CrossClockStdLogic of CrossClockStdLogic is
begin


end behavioral_CrossClockStdLogic;

